* NGSPICE file created from user_proj_example.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180_sram_8x1024 abstract view
.subckt gf180_sram_8x1024 csb0 web0 clk0 dout0[7] addr0[4] addr0[5] addr0[6] addr0[7]
+ addr0[8] addr0[9] vdd gnd din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6]
+ din0[7] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] addr0[0]
+ addr0[1] addr0[2] addr0[3]
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4]
+ io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[1] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[2] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] vdd vss io_out[17] io_out[16]
+ io_out[15] io_out[14] io_oeb[27] io_out[13] io_oeb[26] io_out[12] io_oeb[25] io_out[11]
+ io_oeb[24] io_out[21] io_out[10] irq[2] io_oeb[23] io_out[20] io_oeb[12] irq[1]
+ io_oeb[22] io_out[19] io_oeb[11] irq[0] io_oeb[21] io_out[18] io_oeb[10] io_oeb[20]
+ io_oeb[28]
XFILLER_0_39_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_2_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_187_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_49_2_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_196_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_137_2_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_1_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_1_Right_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_167_1_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_1_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_1_Right_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_127_1_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_2_Left_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_59_1_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_188_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_173_1_Left_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_141_2_Left_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_2_Left_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_1_Right_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_2_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_152_2_Right_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_din0[7] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_2_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_2_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_185_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_1_Right_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_2_Right_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_150_2_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_136_1_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_185_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_1_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_1_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_68_1_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_36_2_Left_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_150_2_Left_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_65_1_Right_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_154_2_Right_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_31_2_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_82_2_Left_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_2_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_2_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_112_2_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_2_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_66_1_Right_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_155_2_Right_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_1_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_2_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_1_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_1_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_1_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_145_1_Left_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_1_Right_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_156_2_Right_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_173_1_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_108_2_Left_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_2_Left_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_77_1_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_194_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_188_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_91_2_Left_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_185_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_191_Left_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_54_1_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_157_2_Right_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_2_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_2_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_din0[6] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_1_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_2_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_108_1_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_158_2_Right_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_1_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_154_1_Left_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_122_2_Left_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_150_2_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_117_2_Left_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_86_1_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_1_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_2_Left_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_180_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_158_1_Right_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_159_2_Right_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_2_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_120_1_Right_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I io_in[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_1_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_2_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_174_2_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_159_1_Right_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input3_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_117_1_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_121_1_Right_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_1_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_1_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_2_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_131_2_Left_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_143_2_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_163_1_Left_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_1_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_63_2_Left_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_95_1_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_85_1_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_173_1_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_122_1_Right_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_2_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_2_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_123_1_Right_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_din0[5] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_2_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_126_1_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_2_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_2_Left_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_58_1_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_172_1_Left_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_140_2_Left_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_185_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_124_1_Right_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_1_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_72_2_Left_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_101_2_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_2_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_125_1_Right_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_1_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_1_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput22 net22 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_198_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_135_1_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_126_1_Right_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_125_2_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_1_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_2_Left_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_88_1_Right_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_183_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_81_2_Left_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_1_Right_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_127_1_Right_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_2_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_2_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_1_Right_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_188_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_51_1_Right_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_din0[4] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_144_1_Left_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_2_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_2_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_2_Left_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_2_Left_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_76_1_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_173_2_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_1_Right_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_148_1_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_2_Left_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_185_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_50_1_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_188_Left_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_53_1_Right_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_197_Left_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_1_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_1_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_2_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_39_1_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput23 net23 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_54_1_Right_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_132_2_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_1_Left_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_121_2_Left_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_2_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_116_2_Left_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_85_1_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_53_2_Left_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_1_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_2_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_192_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_55_1_Right_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_2_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_181_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_1_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_56_1_Right_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_91_1_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_116_1_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_2_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_1_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_100_1_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_130_2_Left_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_162_1_Left_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_1_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_din0[3] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_2_Left_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_94_1_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_1_Right_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_2_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_2_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_148_1_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_1_Right_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_140_2_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_29_1_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_179_1_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_gf180_sram_8x1024_web0 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_2_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_125_1_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_2_Left_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_1_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_2_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_141_2_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput24 net24 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_198_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_71_2_Left_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_103_2_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_162_1_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_32_2_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_148_1_Right_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_192_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_104_2_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_156_2_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_181_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_194_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_149_1_Right_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_134_1_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_190_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_1_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_34_2_Left_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_2_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_2_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_198_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_80_2_Left_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_gf180_sram_8x1024_din0[2] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_106_2_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_1_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_143_1_Left_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_179_1_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_2_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_2_Left_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_2_Left_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_75_1_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput25 net25 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_198_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_108_2_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_2_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_1_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_80_1_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_106_1_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_109_2_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_1_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_1_Right_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_152_1_Left_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_120_2_Left_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_2_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_194_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_115_2_Left_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_84_1_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_2_Left_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_107_2_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_162_2_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_1_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_198_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_71_1_Right_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_183_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_din0[1] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_2_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_72_1_Right_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_1_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_185_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_1_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_1_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_2_Left_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_1_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_2_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_73_1_Right_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_162_2_Right_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_1_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_184_Left_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_193_Left_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_1_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_2_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput26 net26 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_195_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_74_1_Right_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_197_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_163_2_Right_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_145_2_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_2_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_1_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_124_1_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_175_1_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_1400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_24_2_Left_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_1_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_75_1_Right_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_164_2_Right_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_2_Left_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_2_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_2_Left_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_2_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_2_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_162_2_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_1_Right_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_165_2_Right_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_1_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output26_I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_din0[0] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_138_2_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_2_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_19_1_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_77_1_Right_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_168_1_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_166_2_Right_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_1_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_189_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_65_1_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_2_Left_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_167_2_Right_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_2_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_1_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_1_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput27 net27 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_168_2_Right_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_28_1_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_192_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_2_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_142_1_Left_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_105_2_Left_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_2_Left_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_74_1_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_175_1_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_168_1_Right_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_169_2_Right_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_1_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_1_Right_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_81_2_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_130_1_Right_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_194_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_169_1_Right_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_2_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_113_2_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_131_1_Right_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_105_1_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_80 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_187_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_37_1_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_1_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_2_Left_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_83_1_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_2_Left_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_1_Right_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_189_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_1_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input18_I io_in[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_1_Right_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_2_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_2_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_114_1_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput28 net28 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_99_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_1_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_98_2_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_134_1_Right_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_60_2_Left_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_92_1_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_90_2_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_192_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_192_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_1_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_135_1_Right_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_91_2_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_2_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_81_2_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_1_Right_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_2_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_123_1_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_198_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_2_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_98_1_Right_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_23_2_Left_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_55_1_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_70 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_187_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_81 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_138_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_2_Left_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_143_1_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_2_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_137_1_Right_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_99_1_Right_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_1_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_174_1_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_186_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_195_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_2_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_194_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_1_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_168_2_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_1_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_2_Left_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput29 net29 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_2_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_1_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_clk0 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_2_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_181_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_2_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_2_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_1_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_157_1_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_62_1_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_104_2_Left_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_41_2_Left_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_73_1_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_198_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_175_2_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_60 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_71 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_187_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_82 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_198_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_56_2_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_174_1_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_104_1_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_28_1_Right_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_2_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_1_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_2_Left_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_1_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_50_2_Left_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_168_2_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_29_1_Right_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_1_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_150_2_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_2_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_192_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_181_Left_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_112_2_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_190_Left_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_192_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_113_1_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_102_2_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_1_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_2_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_151_2_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_185_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_181_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_1_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_178_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_2_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_157_1_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_61 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_50 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_72 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_138_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_114_2_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_2_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_182_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_189_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_122_1_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_2_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_37_1_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_2_Left_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_1_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_2_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_1_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_116_2_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input16_I io_in[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_1_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_1_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_1_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_117_2_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_63_1_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_102_2_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_2_Left_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_2_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_1_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_194_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_118_2_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_2_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_108_1_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_62 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_51 irq[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_103_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_40 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_73 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_74_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_1_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_119_2_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_80_1_Right_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_1_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_189_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_2_Left_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_40_2_Left_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_72_1_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_157_2_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_1_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_81_1_Right_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_179_2_Left_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_1_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput1 io_in[10] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_174_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_2_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_61_2_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_1_Right_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_103_1_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_170_1_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_1_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_1_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_1_Right_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_112_2_Left_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_2_Right_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_1_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_2_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_2_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_84_1_Right_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_173_2_Right_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_2_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_70_2_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_30 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_52 irq[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_75_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_41 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_63 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_74 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_187_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_163_1_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_112_1_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_1_Right_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_187_Left_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_44_1_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_174_2_Right_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_196_Left_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_189_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_2_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_2_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_86_1_Right_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_175_2_Right_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput2 io_in[11] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_8_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_2_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_1_Right_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_68_1_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_176_2_Right_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_185_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_2_Left_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_1_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_121_1_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_177_2_Right_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_196_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input21_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_192_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_2_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_178_2_Right_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_2_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_31 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_53 irq[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_42 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_177_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_64 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_75 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_198_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_51_2_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_62_1_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_2_Left_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_178_1_Right_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_179_2_Right_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_6_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_169_2_Left_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_140_1_Right_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_182_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_188_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_179_1_Right_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_2_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_141_1_Right_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 io_in[12] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_163_2_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_1_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_1_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_102_2_Left_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_142_1_Right_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_1_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_178_2_Left_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_1_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_196_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_143_1_Right_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input14_I io_in[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_2_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_60_2_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_152_1_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_185_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_102_1_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_2_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_144_1_Right_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_1_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_1_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_111_2_Left_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_example_32 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_100_2_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_43 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_65 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_54 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_76 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_187_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_146_2_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_2_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_addr0[9] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_145_1_Right_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_1_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_182_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_2_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_2_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_146_1_Right_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_2_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 io_in[13] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_163_2_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_108_1_Right_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_1_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_1_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_147_1_Right_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_171_1_Left_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_19_1_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_109_1_Right_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_169_1_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_196_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_34_2_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_152_1_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_185_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_20_2_Left_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_1_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_98_1_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_159_2_Left_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_180_1_Left_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_33 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_44 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_66 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_77 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_55 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_2_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_6_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_189_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_gf180_sram_8x1024_addr0[8] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_197_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_2_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_198_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_176_1_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_182_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_188_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_1_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_183_Left_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_2_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_192_Left_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[14] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_2_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_168_2_Left_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_110_1_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_1_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_169_1_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_2_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_1_Right_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_1_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_129_2_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_2_Left_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_191_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_2_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_1_Right_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_177_2_Left_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_103_1_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_193_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_160_2_Right_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_34 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_103_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_78 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_45 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_56 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_187_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_67 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_74_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_6_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_2_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_gf180_sram_8x1024_addr0[7] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_197_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_2_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_1_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_1_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_160_1_Right_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_161_2_Right_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_1_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_110_2_Left_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_123_2_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_161_1_Left_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_2_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput6 io_in[15] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_161_1_Right_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_26_2_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_2_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_1_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_124_2_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_1_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_2_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_1_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_162_1_Right_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_2_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_104_2_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_2_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_1_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_42_1_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput20 io_in[8] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_149_2_Left_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_163_1_Right_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_170_1_Left_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_2_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_2_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_126_2_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_103_1_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_1_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I io_in[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_2_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_164_1_Right_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_35 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_46 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_57 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_68 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_input4_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_79 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_146_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_127_2_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_146_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_addr0[6] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_2_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_165_1_Right_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_182_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_1_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_158_2_Left_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_128_2_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_2_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_166_1_Right_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput7 io_in[16] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_38_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_1_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_40_2_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_129_2_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_176_2_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_1_Right_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_167_1_Right_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_1_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_2_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_87_1_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_1_Right_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_196_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput21 io_in[9] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput10 io_in[19] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_167_2_Left_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_110_2_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_2_Left_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_191_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_191_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_1_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_2_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_1_Left_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_92_1_Right_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_1_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_1_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_23_1_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_36 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_47 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_69 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_58 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_177_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_6_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_93_1_Right_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_100_2_Left_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_addr0[5] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_1_Left_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_197_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_2_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_176_2_Left_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_185_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_194_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_2_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_1_Right_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_1_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_1_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_2_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[17] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_188_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_158_1_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_95_1_Right_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_1_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_2_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_139_2_Left_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_160_1_Left_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_96_1_Right_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput11 io_in[20] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_1_Right_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_2_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_1_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_93_1_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_88_2_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_2_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_1_Right_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_97_1_Right_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_140_1_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_59_1_Right_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_1_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_1_Right_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_171_1_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_example_59 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_37 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_48 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_148_2_Left_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_addr0[4] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_186_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_182_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_1_Right_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_30_2_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_2_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_2_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_2_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_1_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_133_1_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_in[18] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_160_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_23_1_Right_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_2_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_1_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_76_1_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_1_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_150_1_Right_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_127_2_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_157_2_Left_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_1_Right_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_89_2_Left_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_1_Right_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_196_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_2_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput12 io_in[21] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_1_Right_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_189_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_152_1_Right_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_1_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_1_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_141_2_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_1_Right_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_166_2_Left_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_184_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_1_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_example_49 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_38 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_190_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_98_2_Left_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_2_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_153_1_Right_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_gf180_sram_8x1024_addr0[3] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_84_2_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input10_I io_in[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_59_2_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_1_Right_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_186_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_52_1_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input2_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_165_2_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_154_1_Right_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_1_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_2_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_110_2_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_129_2_Left_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_2_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_150_1_Left_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_109_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_155_1_Right_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_175_2_Left_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_1_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_164_1_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_194_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_111_2_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_179_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_68_2_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_156_1_Right_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_158_2_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput13 io_in[22] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_1_Right_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_191_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_157_1_Right_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_1_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_138_2_Left_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_189_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_10_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_1_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_1_Right_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_2_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_proj_example_39 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_197_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_2_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_77_2_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_addr0[2] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_179_2_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_2_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_2_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_186_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_2_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_179_1_Left_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_147_2_Left_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_2_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_79_2_Left_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_146_1_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_2_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_27_1_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput14 io_in[23] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_184_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_131_1_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_2_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_2_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_156_2_Left_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_1_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_191_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_1_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_2_Left_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_189_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_186_Left_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_195_Left_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_49_2_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_48_1_Right_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_2_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_1_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_addr0[1] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_2_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_186_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_2_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_140_1_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_1_Right_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_90_2_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_165_2_Left_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_153_1_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_2_Left_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_2_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_170_2_Right_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_2_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_2_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_2_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_2_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_2_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_182_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_191_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_1_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_170_1_Right_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_171_2_Right_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_177_1_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_2_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_128_2_Left_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput15 io_in[24] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_58_1_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_81_1_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_171_1_Right_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_130_2_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_174_2_Left_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_160_1_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_195_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_2_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_195_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_191_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_1_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_67_2_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_1_Right_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_184_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_135_2_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_gf180_sram_8x1024_addr0[0] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_197_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_173_1_Right_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_137_2_Left_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_169_1_Left_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_2_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_2_Left_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_90_1_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_136_2_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_153_1_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_174_1_Right_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_1_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_76_2_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_2_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_122_2_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_2_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_2_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_175_1_Right_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_121_1_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_1_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_138_2_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_178_1_Left_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_146_2_Left_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_2_Left_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_2_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_176_1_Right_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput16 io_in[25] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_58_1_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_2_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_139_2_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I io_in[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_2_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_100_1_Right_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_111_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_177_1_Right_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_130_1_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_101_1_Right_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_155_2_Left_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_197_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_87_2_Left_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_1_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_17_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_48_2_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_102_1_Right_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_2_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_122_2_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_1_Right_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_1_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_164_2_Left_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_2_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_2_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_96_2_Left_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_179_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_104_1_Right_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_1_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_csb0 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_2_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput17 io_in[26] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_105_1_Right_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_195_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_191_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_2_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_189_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_177_2_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_188_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_197_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_159_1_Left_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_127_2_Left_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_185_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_184_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_59_2_Left_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_182_Left_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_192_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_1_Right_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_1_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_173_2_Left_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_2_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_68_1_Right_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_105_2_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_88_1_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_30_1_Right_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_2_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_135_1_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_107_1_Right_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_146_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_69_1_Right_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_41_2_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_31_1_Right_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_104_1_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_111_1_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_1_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_136_2_Left_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_168_1_Left_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_68_2_Left_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_1_Right_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_2_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_2_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_1_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_75_2_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_95_1_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output25_I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput18 io_in[27] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_1_Right_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_120_1_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_195_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_1_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_1773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_2_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_177_1_Left_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_145_2_Left_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_1_Right_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_77_2_Left_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_184_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_38_2_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_58_2_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_35_1_Right_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_88_1_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_141_1_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_36_1_Right_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_61_1_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_2_Left_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_1_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_dout0[7] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xgf180_sram_8x1024 net18 net17 net19 net29 net11 net12 net13 net14 net15 net16 vdd
+ vss net20 net21 net1 net2 net3 net4 net5 net6 net22 net23 net24 net25 net26 net27
+ net28 net7 net8 net9 net10 gf180_sram_8x1024
XFILLER_0_113_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_86_2_Left_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_1_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_2_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_37_1_Right_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_2_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput19 io_in[28] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_120_2_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_1_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_1_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_149_1_Left_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_2_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_49_2_Left_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_70_1_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_159_1_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_163_2_Left_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_2_Left_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_121_2_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_83_2_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_56_2_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input17_I io_in[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_2_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_128_1_Right_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I io_in[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_84_2_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_1_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_186_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_158_1_Left_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_126_2_Left_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_129_1_Right_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_1_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_2_Left_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_2_Left_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_2_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_2_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_gf180_sram_8x1024_dout0[6] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_2_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_1_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_65_2_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_1_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_86_2_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_1_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_110_1_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_166_2_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_135_2_Left_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_167_1_Left_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_2_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_1_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_67_2_Left_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_99_1_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_185_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_2_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_2_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_1_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_88_2_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_74_2_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_184_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_184_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_193_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_30_2_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_2_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_2_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_1_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_51_1_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_60_1_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_5_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_176_1_Left_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_186_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_144_2_Left_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_1_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_2_Left_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_2_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_2_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_2_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_dout0[5] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_142_2_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_1_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_172_1_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_1_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_189_Left_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_39_2_Left_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_1_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_198_Left_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_1_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_153_2_Left_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_2_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_85_2_Left_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_180_2_Right_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_2_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_142_2_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_46_2_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_195_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_2_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output23_I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_180_1_Right_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_1_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_190_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_190_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_143_2_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_148_1_Left_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_1_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_2_Left_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_180_2_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_162_2_Left_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_1_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_5_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_144_2_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_186_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_2_Left_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_55_2_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_145_2_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_149_2_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_gf180_sram_8x1024_dout0[4] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_2_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_157_1_Left_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_125_2_Left_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_123_1_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_146_2_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_89_1_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_2_Left_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_171_2_Left_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_18_2_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_64_2_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_117_2_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_2_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_147_2_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_147_1_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_3_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_2_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_148_2_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_190_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_190_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_41_1_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_1_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_134_2_Left_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_166_1_Left_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_66_2_Left_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_98_1_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_180_2_Left_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_130_1_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_2_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_149_2_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_131_2_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input15_I io_in[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_2_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_110_1_Right_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_77_2_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_1_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_124_2_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I io_in[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_gf180_sram_8x1024_dout0[3] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_129_1_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_111_1_Right_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_2_Left_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_1_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_175_1_Left_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_143_2_Left_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_155_2_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_2_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_75_2_Left_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_1_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_112_1_Right_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_2_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_2_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_1_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_1_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_2_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_1_Right_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_1_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_138_1_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_38_2_Left_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_152_2_Left_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_2_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_190_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_1_Right_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_84_2_Left_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_1_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_45_2_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_1_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_115_1_Right_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_131_2_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_77_2_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_1_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_179_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_181_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_147_1_Left_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_116_1_Right_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_gf180_sram_8x1024_dout0[2] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_2_Left_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_79_1_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_161_2_Left_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_78_1_Right_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_2_Left_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_2_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_1_Right_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_54_2_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_117_1_Right_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_79_1_Right_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_1_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_2_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_91_2_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_41_1_Right_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_185_Left_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_1_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_194_Left_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_31_1_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_156_1_Left_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_124_2_Left_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_195_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_195_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_2_Left_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_88_1_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_56_2_Left_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_2_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_170_2_Left_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_42_1_Right_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_148_2_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_190_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_178_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_63_2_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_1_Right_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_1_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_119_1_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_1_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_44_1_Right_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_2_Left_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_165_1_Left_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_2_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_181_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_181_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_2_Left_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_97_1_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_190_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input20_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_gf180_sram_8x1024_dout0[1] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_2_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_45_1_Right_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_72_2_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_174_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_194_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_2_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_1_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_46_1_Right_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_128_1_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_193_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_28_2_Left_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_2_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_195_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_174_1_Left_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_142_2_Left_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_74_2_Left_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_47_1_Right_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_2_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_2_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_188_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_1_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_130_2_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_1_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_1_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_92_2_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_137_1_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_183_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_1_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_37_2_Left_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_151_2_Left_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_131_2_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_2_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_83_2_Left_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_2_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_93_2_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_44_2_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_gf180_sram_8x1024_dout0[0] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input13_I io_in[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_1_Right_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_2_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input5_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_94_2_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_106_2_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_2_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_1_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_146_1_Left_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_1650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_1_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_1_Right_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_172_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_109_2_Left_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_2_Left_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_78_1_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_160_2_Left_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_95_2_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_2_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_2_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_2_Left_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_167_1_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_195_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_2_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_190_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_2_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_1_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_150_1_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_1_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_155_1_Left_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_198_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_2_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_123_2_Left_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_1_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_2_Left_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_183_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_1_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_183_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_55_2_Left_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_2_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_2_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_178_2_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_2_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_118_1_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_1_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_198_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_1_Right_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_132_2_Left_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_164_1_Left_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_1_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_2_Left_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_96_1_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_24_2_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

