VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1030.660 BY 800.320 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 28.000 1030.660 28.560 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 796.320 552.720 800.320 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 796.320 438.480 800.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 796.320 324.240 800.320 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 796.320 210.000 800.320 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 796.320 95.760 800.320 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 789.600 4.000 790.160 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 732.480 4.000 733.040 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.360 4.000 675.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.240 4.000 618.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 159.040 1030.660 159.600 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 4.000 447.440 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.760 4.000 390.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END io_in[28]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 290.080 1030.660 290.640 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 421.120 1030.660 421.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 552.160 1030.660 552.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 683.200 1030.660 683.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1009.120 796.320 1009.680 800.320 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.880 796.320 895.440 800.320 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 796.320 781.200 800.320 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 796.320 666.960 800.320 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 115.360 1030.660 115.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 796.320 476.560 800.320 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 796.320 362.320 800.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 796.320 248.080 800.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 796.320 133.840 800.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 796.320 19.600 800.320 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 751.520 4.000 752.080 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.280 4.000 637.840 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 580.160 4.000 580.720 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 523.040 4.000 523.600 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 246.400 1030.660 246.960 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 465.920 4.000 466.480 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.680 4.000 352.240 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.560 4.000 295.120 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.440 4.000 238.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.960 4.000 9.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 377.440 1030.660 378.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 508.480 1030.660 509.040 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 639.520 1030.660 640.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 770.560 1030.660 771.120 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 932.960 796.320 933.520 800.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 818.720 796.320 819.280 800.320 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 796.320 705.040 800.320 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 796.320 590.800 800.320 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 71.680 1030.660 72.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 796.320 514.640 800.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 796.320 400.400 800.320 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 796.320 286.160 800.320 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 796.320 171.920 800.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 796.320 57.680 800.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.560 4.000 771.120 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 713.440 4.000 714.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 656.320 4.000 656.880 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 599.200 4.000 599.760 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 542.080 4.000 542.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 202.720 1030.660 203.280 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.960 4.000 485.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 427.840 4.000 428.400 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 370.720 4.000 371.280 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 4.000 28.560 ;
    END
  END io_out[28]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 333.760 1030.660 334.320 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 464.800 1030.660 465.360 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 595.840 1030.660 596.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1026.660 726.880 1030.660 727.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 796.320 971.600 800.320 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 796.320 857.360 800.320 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 796.320 743.120 800.320 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 796.320 628.880 800.320 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 0.000 514.640 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 0.000 857.360 4.000 ;
    END
  END irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 100.325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 714.775 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 89.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 199.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 105.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 176.920 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 25.540 15.380 27.140 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 15.380 180.740 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 15.380 334.340 100.325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 176.920 334.340 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 15.380 487.940 105.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 176.920 487.940 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.940 15.380 641.540 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 793.540 15.380 795.140 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 947.140 15.380 948.740 784.300 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1023.680 787.210 ;
      LAYER Metal2 ;
        RECT 8.540 796.020 18.740 796.320 ;
        RECT 19.900 796.020 56.820 796.320 ;
        RECT 57.980 796.020 94.900 796.320 ;
        RECT 96.060 796.020 132.980 796.320 ;
        RECT 134.140 796.020 171.060 796.320 ;
        RECT 172.220 796.020 209.140 796.320 ;
        RECT 210.300 796.020 247.220 796.320 ;
        RECT 248.380 796.020 285.300 796.320 ;
        RECT 286.460 796.020 323.380 796.320 ;
        RECT 324.540 796.020 361.460 796.320 ;
        RECT 362.620 796.020 399.540 796.320 ;
        RECT 400.700 796.020 437.620 796.320 ;
        RECT 438.780 796.020 475.700 796.320 ;
        RECT 476.860 796.020 513.780 796.320 ;
        RECT 514.940 796.020 551.860 796.320 ;
        RECT 553.020 796.020 589.940 796.320 ;
        RECT 591.100 796.020 628.020 796.320 ;
        RECT 629.180 796.020 666.100 796.320 ;
        RECT 667.260 796.020 704.180 796.320 ;
        RECT 705.340 796.020 742.260 796.320 ;
        RECT 743.420 796.020 780.340 796.320 ;
        RECT 781.500 796.020 818.420 796.320 ;
        RECT 819.580 796.020 856.500 796.320 ;
        RECT 857.660 796.020 894.580 796.320 ;
        RECT 895.740 796.020 932.660 796.320 ;
        RECT 933.820 796.020 970.740 796.320 ;
        RECT 971.900 796.020 1008.820 796.320 ;
        RECT 1009.980 796.020 1021.860 796.320 ;
        RECT 8.540 4.300 1021.860 796.020 ;
        RECT 8.540 4.000 171.060 4.300 ;
        RECT 172.220 4.000 513.780 4.300 ;
        RECT 514.940 4.000 856.500 4.300 ;
        RECT 857.660 4.000 1021.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 789.300 1026.660 790.020 ;
        RECT 4.000 771.420 1026.660 789.300 ;
        RECT 4.300 770.260 1026.360 771.420 ;
        RECT 4.000 752.380 1026.660 770.260 ;
        RECT 4.300 751.220 1026.660 752.380 ;
        RECT 4.000 733.340 1026.660 751.220 ;
        RECT 4.300 732.180 1026.660 733.340 ;
        RECT 4.000 727.740 1026.660 732.180 ;
        RECT 4.000 726.580 1026.360 727.740 ;
        RECT 4.000 714.300 1026.660 726.580 ;
        RECT 4.300 713.140 1026.660 714.300 ;
        RECT 4.000 695.260 1026.660 713.140 ;
        RECT 4.300 694.100 1026.660 695.260 ;
        RECT 4.000 684.060 1026.660 694.100 ;
        RECT 4.000 682.900 1026.360 684.060 ;
        RECT 4.000 676.220 1026.660 682.900 ;
        RECT 4.300 675.060 1026.660 676.220 ;
        RECT 4.000 657.180 1026.660 675.060 ;
        RECT 4.300 656.020 1026.660 657.180 ;
        RECT 4.000 640.380 1026.660 656.020 ;
        RECT 4.000 639.220 1026.360 640.380 ;
        RECT 4.000 638.140 1026.660 639.220 ;
        RECT 4.300 636.980 1026.660 638.140 ;
        RECT 4.000 619.100 1026.660 636.980 ;
        RECT 4.300 617.940 1026.660 619.100 ;
        RECT 4.000 600.060 1026.660 617.940 ;
        RECT 4.300 598.900 1026.660 600.060 ;
        RECT 4.000 596.700 1026.660 598.900 ;
        RECT 4.000 595.540 1026.360 596.700 ;
        RECT 4.000 581.020 1026.660 595.540 ;
        RECT 4.300 579.860 1026.660 581.020 ;
        RECT 4.000 561.980 1026.660 579.860 ;
        RECT 4.300 560.820 1026.660 561.980 ;
        RECT 4.000 553.020 1026.660 560.820 ;
        RECT 4.000 551.860 1026.360 553.020 ;
        RECT 4.000 542.940 1026.660 551.860 ;
        RECT 4.300 541.780 1026.660 542.940 ;
        RECT 4.000 523.900 1026.660 541.780 ;
        RECT 4.300 522.740 1026.660 523.900 ;
        RECT 4.000 509.340 1026.660 522.740 ;
        RECT 4.000 508.180 1026.360 509.340 ;
        RECT 4.000 504.860 1026.660 508.180 ;
        RECT 4.300 503.700 1026.660 504.860 ;
        RECT 4.000 485.820 1026.660 503.700 ;
        RECT 4.300 484.660 1026.660 485.820 ;
        RECT 4.000 466.780 1026.660 484.660 ;
        RECT 4.300 465.660 1026.660 466.780 ;
        RECT 4.300 465.620 1026.360 465.660 ;
        RECT 4.000 464.500 1026.360 465.620 ;
        RECT 4.000 447.740 1026.660 464.500 ;
        RECT 4.300 446.580 1026.660 447.740 ;
        RECT 4.000 428.700 1026.660 446.580 ;
        RECT 4.300 427.540 1026.660 428.700 ;
        RECT 4.000 421.980 1026.660 427.540 ;
        RECT 4.000 420.820 1026.360 421.980 ;
        RECT 4.000 409.660 1026.660 420.820 ;
        RECT 4.300 408.500 1026.660 409.660 ;
        RECT 4.000 390.620 1026.660 408.500 ;
        RECT 4.300 389.460 1026.660 390.620 ;
        RECT 4.000 378.300 1026.660 389.460 ;
        RECT 4.000 377.140 1026.360 378.300 ;
        RECT 4.000 371.580 1026.660 377.140 ;
        RECT 4.300 370.420 1026.660 371.580 ;
        RECT 4.000 352.540 1026.660 370.420 ;
        RECT 4.300 351.380 1026.660 352.540 ;
        RECT 4.000 334.620 1026.660 351.380 ;
        RECT 4.000 333.500 1026.360 334.620 ;
        RECT 4.300 333.460 1026.360 333.500 ;
        RECT 4.300 332.340 1026.660 333.460 ;
        RECT 4.000 314.460 1026.660 332.340 ;
        RECT 4.300 313.300 1026.660 314.460 ;
        RECT 4.000 295.420 1026.660 313.300 ;
        RECT 4.300 294.260 1026.660 295.420 ;
        RECT 4.000 290.940 1026.660 294.260 ;
        RECT 4.000 289.780 1026.360 290.940 ;
        RECT 4.000 276.380 1026.660 289.780 ;
        RECT 4.300 275.220 1026.660 276.380 ;
        RECT 4.000 257.340 1026.660 275.220 ;
        RECT 4.300 256.180 1026.660 257.340 ;
        RECT 4.000 247.260 1026.660 256.180 ;
        RECT 4.000 246.100 1026.360 247.260 ;
        RECT 4.000 238.300 1026.660 246.100 ;
        RECT 4.300 237.140 1026.660 238.300 ;
        RECT 4.000 219.260 1026.660 237.140 ;
        RECT 4.300 218.100 1026.660 219.260 ;
        RECT 4.000 203.580 1026.660 218.100 ;
        RECT 4.000 202.420 1026.360 203.580 ;
        RECT 4.000 200.220 1026.660 202.420 ;
        RECT 4.300 199.060 1026.660 200.220 ;
        RECT 4.000 181.180 1026.660 199.060 ;
        RECT 4.300 180.020 1026.660 181.180 ;
        RECT 4.000 162.140 1026.660 180.020 ;
        RECT 4.300 160.980 1026.660 162.140 ;
        RECT 4.000 159.900 1026.660 160.980 ;
        RECT 4.000 158.740 1026.360 159.900 ;
        RECT 4.000 143.100 1026.660 158.740 ;
        RECT 4.300 141.940 1026.660 143.100 ;
        RECT 4.000 124.060 1026.660 141.940 ;
        RECT 4.300 122.900 1026.660 124.060 ;
        RECT 4.000 116.220 1026.660 122.900 ;
        RECT 4.000 115.060 1026.360 116.220 ;
        RECT 4.000 105.020 1026.660 115.060 ;
        RECT 4.300 103.860 1026.660 105.020 ;
        RECT 4.000 85.980 1026.660 103.860 ;
        RECT 4.300 84.820 1026.660 85.980 ;
        RECT 4.000 72.540 1026.660 84.820 ;
        RECT 4.000 71.380 1026.360 72.540 ;
        RECT 4.000 66.940 1026.660 71.380 ;
        RECT 4.300 65.780 1026.660 66.940 ;
        RECT 4.000 47.900 1026.660 65.780 ;
        RECT 4.300 46.740 1026.660 47.900 ;
        RECT 4.000 28.860 1026.660 46.740 ;
        RECT 4.300 27.700 1026.360 28.860 ;
        RECT 4.000 9.820 1026.660 27.700 ;
        RECT 4.300 9.100 1026.660 9.820 ;
      LAYER Metal4 ;
        RECT 100.000 84.090 175.540 712.860 ;
        RECT 177.740 84.090 178.840 712.860 ;
        RECT 181.040 176.620 332.440 712.860 ;
        RECT 334.640 199.080 482.740 712.860 ;
        RECT 484.940 199.080 486.040 712.860 ;
        RECT 334.640 176.620 486.040 199.080 ;
        RECT 488.240 176.620 636.340 712.860 ;
        RECT 638.540 176.620 639.640 712.860 ;
        RECT 181.040 106.240 639.640 176.620 ;
        RECT 181.040 105.580 636.340 106.240 ;
        RECT 181.040 100.625 486.040 105.580 ;
        RECT 181.040 84.090 329.140 100.625 ;
        RECT 331.340 84.090 332.440 100.625 ;
        RECT 334.640 89.740 486.040 100.625 ;
        RECT 334.640 84.090 482.740 89.740 ;
        RECT 484.940 84.090 486.040 89.740 ;
        RECT 488.240 84.090 636.340 105.580 ;
        RECT 638.540 84.090 639.640 106.240 ;
        RECT 641.840 84.090 789.940 712.860 ;
        RECT 792.140 84.090 793.240 712.860 ;
        RECT 795.440 84.090 931.320 712.860 ;
  END
END user_proj_example
END LIBRARY

