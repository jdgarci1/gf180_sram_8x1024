// This is the unpowered netlist.
module user_proj_example (io_in,
    io_oeb,
    io_out,
    irq);
 input [28:0] io_in;
 output [28:0] io_oeb;
 output [28:0] io_out;
 output [2:0] irq;

 wire net54;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net55;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net81;
 wire net82;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net30;
 wire net31;
 wire net51;
 wire net52;
 wire net53;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[0]  (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[1]  (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[2]  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[3]  (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[4]  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[5]  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[6]  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[7]  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[8]  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_addr0[9]  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf180_sram_8x1024_clk0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf180_sram_8x1024_csb0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[0]  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[1]  (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[2]  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[3]  (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[4]  (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[5]  (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[6]  (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_din0[7]  (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[0]  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[1]  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[2]  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[3]  (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[4]  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[5]  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[6]  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_gf180_sram_8x1024_dout0[7]  (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_gf180_sram_8x1024_web0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_183_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_183_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_184_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_184_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_185_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_185_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_185_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_185_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_186_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_187_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_187_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_187_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_188_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_188_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_189_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_189_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_189_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_189_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_190_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_190_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_191_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_191_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_191_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_191_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_192_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_195_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_196_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_196_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_196_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_197_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_197_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_197_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_197_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_197_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_198_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_198_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_198_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_198_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_1_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_1_Right_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Left_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_2_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_1_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_1_Right_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Left_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_2_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_1_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_1_Right_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Left_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_2_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_1_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_1_Right_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Left_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_2_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_1_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_1_Right_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Left_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_2_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_1_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_1_Right_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Left_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_2_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_1_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_1_Right_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Left_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_2_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_1_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_1_Right_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Left_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_2_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_1_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_1_Right_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Left_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_2_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_1_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_1_Right_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Left_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_2_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_1_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_1_Right_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Left_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_2_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_1_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_1_Right_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Left_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_2_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_1_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_1_Right_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Left_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_2_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_1_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_1_Right_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Left_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_2_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_1_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_1_Right_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Left_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_2_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_1_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_1_Right_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Left_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_2_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_1_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_1_Right_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Left_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_2_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_1_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_1_Right_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Left_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_2_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_1_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_1_Right_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Left_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_2_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_1_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_1_Right_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Left_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_2_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_1_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_1_Right_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Left_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_2_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_1_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_1_Right_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Left_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_2_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_1_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_1_Right_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Left_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_2_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_1_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_1_Right_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Left_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_2_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_1_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_1_Right_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Left_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_2_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_1_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_1_Right_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Left_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_2_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_1_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_1_Right_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Left_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_2_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_1_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_1_Right_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Left_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_2_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_1_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_1_Right_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Left_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_2_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_1_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_1_Right_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Left_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_2_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_1_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_1_Right_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Left_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_2_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_1_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_1_Right_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Left_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_2_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_1_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_1_Right_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Left_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_2_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_1_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_1_Right_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Left_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_2_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_1_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_1_Right_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Left_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_2_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_1_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_1_Right_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Left_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_2_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_1_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_1_Right_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Left_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_2_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_1_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_1_Right_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Left_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_2_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_1_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_1_Right_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Left_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_2_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_1_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_1_Right_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Left_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_2_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_1_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_1_Right_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Left_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_2_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_1_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_1_Right_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Left_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_2_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_1_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_1_Right_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Left_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_2_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_1_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_1_Right_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Left_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_2_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_1_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_1_Right_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Left_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_2_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_1_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_1_Right_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Left_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_2_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_1_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_1_Right_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Left_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_2_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_1_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_1_Right_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Left_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_2_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_1_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_1_Right_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Left_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_2_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_1_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_1_Right_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Left_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_2_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_1_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_1_Right_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Left_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_2_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_1_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_1_Right_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Left_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_2_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_1_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_1_Right_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Left_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_2_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_1_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_1_Right_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Left_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_2_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_1_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_1_Right_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Left_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_2_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_1_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_1_Right_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Left_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_2_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_1_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_1_Right_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Left_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_2_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_1_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_1_Right_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Left_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_2_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_1_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_1_Right_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Left_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_2_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_1_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_1_Right_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Left_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_2_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_1_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_1_Right_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Left_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_2_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_1_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_1_Right_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Left_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_2_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_1_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_1_Right_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Left_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_2_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_1_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_1_Right_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Left_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_2_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_1_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_1_Right_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Left_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_2_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_1_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_1_Right_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Left_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_2_Right_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_1_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_1_Right_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Left_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_2_Right_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_1_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_1_Right_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Left_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_2_Right_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_1_Left_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_1_Right_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Left_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_2_Right_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_1_Left_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_1_Right_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Left_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_2_Right_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_1_Left_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_1_Right_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Left_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_2_Right_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_1_Left_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_1_Right_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Left_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_2_Right_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_1_Left_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_1_Right_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Left_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_2_Right_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_1_Left_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_1_Right_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Left_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_2_Right_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_1_Left_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_1_Right_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Left_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_2_Right_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_1_Left_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_1_Right_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Left_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_2_Right_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_1_Left_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_1_Right_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Left_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_2_Right_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_1_Left_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_1_Right_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Left_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_2_Right_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_1_Left_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_1_Right_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Left_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_2_Right_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_1_Left_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_1_Right_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Left_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_2_Right_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_1_Left_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_1_Right_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Left_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_2_Right_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Left_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Left_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Left_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Left_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Left_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Left_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Left_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_1_Left_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_1_Right_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Left_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Left_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Left_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Left_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Left_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Left_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_Left_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_196_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_Left_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_197_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_Left_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_198_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_1_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_1_Right_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_1_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_1_Right_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_1_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_1_Right_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_1_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_1_Right_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_1_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_1_Right_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_1_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_1_Right_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_1_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_1_Right_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_1_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_1_Right_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_1_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_1_Right_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_1_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_1_Right_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_1_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_1_Right_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_1_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_1_Right_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_1_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_1_Right_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_1_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_1_Right_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_1_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_1_Right_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_1_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_1_Right_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_1_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_1_Right_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_1_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_1_Right_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_1_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_1_Right_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_1_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_1_Right_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_1_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_1_Right_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_1_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_1_Right_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_1_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_1_Right_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_1_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_1_Right_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_1_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_1_Right_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_1_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_1_Right_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_1_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_1_Right_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_1_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_1_Right_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_1_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_1_Right_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_1_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_1_Right_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_1_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_1_Right_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_1_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_1_Right_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_1_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_1_Right_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_1_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_1_Right_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_1_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_1_Right_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_1_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_1_Right_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_1_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_1_Right_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_1_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_1_Right_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_1_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_1_Right_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_1_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_1_Right_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_1_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_1_Right_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_1_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_1_Right_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_1_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_1_Right_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_1_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_1_Right_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_1_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_1_Right_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_1_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_1_Right_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_1_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_1_Right_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_1_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_1_Right_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_1_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_1_Right_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_1_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_1_Right_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_1_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_1_Right_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_1_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_1_Right_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_1_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_1_Right_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_1_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_1_Right_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_1_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_1_Right_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_1_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_1_Right_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_1_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_1_Right_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_1_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_1_Right_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_1_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_1_Right_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_1_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_1_Right_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_1_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_1_Right_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_1_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_1_Right_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_1_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_1_Right_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_1_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_1_Right_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_1_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_1_Right_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Left_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_2_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_1_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_1_Right_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Left_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_2_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_1_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_1_Right_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Left_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_2_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_1_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_1_Right_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Left_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_2_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_1_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_1_Right_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Left_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_2_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_1_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_1_Right_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Left_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_2_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_1_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_1_Right_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Left_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_2_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_1_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_1_Right_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Left_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_2_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_1_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_1_Right_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Left_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_2_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_1_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_1_Right_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Left_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_2_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_1_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_1_Right_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Left_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_2_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_1_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_1_Right_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Left_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_2_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_1_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_1_Right_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Left_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_2_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_1_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_1_Right_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Left_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_2_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_1_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_1_Right_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Left_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_2_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_1_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_1_Right_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Left_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_2_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_1_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_1_Right_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Left_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_2_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_1_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_1_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_1_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_1_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_1_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_1_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_1_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_1_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_1_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_1_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_1_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_1_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_1_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_1_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_1_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_1_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_1_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_1_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_1_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_1_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_1_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_1_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_1_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_1_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_1_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_1_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_1_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_1_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_1_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_1_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_1_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_1_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_1_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_1_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_1_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_1_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_1_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_1_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_1_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_1_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_1_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_1_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_1_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_1_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_1_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_1_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_1_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_1_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_1_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_1_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_1_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_1_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_1_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_1_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_1_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_1_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_1_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_1_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_1_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_1_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_1_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_2_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_1_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_1_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_2_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_1_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_1_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_2_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_1_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_1_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_2_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_1_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_1_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_2_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_1_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_1_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_2_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_1_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_1_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_2_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_1_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_1_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_2_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_1_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_1_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_2_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_1_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_1_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_2_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_1_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_1_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_2_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_1_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_2_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_1_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_1_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_2_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_1_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_1_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_2_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_1_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_2_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_1_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_1_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_2_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_1_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_1_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_2_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_1_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_1_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_2_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_1_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_1_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_2_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_1_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_1_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_2_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_1_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_1_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_2_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_1_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_2_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_1_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_1_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_2_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_1_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_2_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_2_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_196_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_197_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_198_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_2_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_2_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_2_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_2_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_2_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_2_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_2_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_2_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_2_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_2_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_2_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_2_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_2_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_2_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_2_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_2_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_2_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_2_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_2_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_2_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_2_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_2_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_2_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_2_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_2_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_2_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_2_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_2_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_2_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_999 ();
 gf180_sram_8x1024 gf180_sram_8x1024 (.csb0(net18),
    .web0(net17),
    .clk0(net19),
    .addr0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9,
    net8,
    net7}),
    .din0({net6,
    net5,
    net4,
    net3,
    net2,
    net1,
    net21,
    net20}),
    .dout0({net29,
    net28,
    net27,
    net26,
    net25,
    net24,
    net23,
    net22}));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input10 (.I(io_in[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(io_in[20]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(io_in[21]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(io_in[22]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(io_in[23]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(io_in[24]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(io_in[25]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(io_in[26]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(io_in[27]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(io_in[28]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input20 (.I(io_in[8]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input21 (.I(io_in[9]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input5 (.I(io_in[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input6 (.I(io_in[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input7 (.I(io_in[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input8 (.I(io_in[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input9 (.I(io_in[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_62 (.Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_63 (.Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_64 (.Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_65 (.Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_66 (.Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_67 (.Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_68 (.Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_69 (.Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_70 (.Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_71 (.Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_72 (.Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_73 (.Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_74 (.Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_75 (.Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_76 (.Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_77 (.Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_78 (.Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_79 (.Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_80 (.Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_81 (.Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_82 (.Z(net82));
 assign io_oeb[0] = net54;
 assign io_oeb[10] = net62;
 assign io_oeb[11] = net63;
 assign io_oeb[12] = net64;
 assign io_oeb[13] = net65;
 assign io_oeb[14] = net66;
 assign io_oeb[15] = net67;
 assign io_oeb[16] = net68;
 assign io_oeb[17] = net69;
 assign io_oeb[18] = net70;
 assign io_oeb[19] = net71;
 assign io_oeb[1] = net55;
 assign io_oeb[20] = net72;
 assign io_oeb[21] = net73;
 assign io_oeb[22] = net74;
 assign io_oeb[23] = net75;
 assign io_oeb[24] = net76;
 assign io_oeb[25] = net77;
 assign io_oeb[26] = net78;
 assign io_oeb[27] = net79;
 assign io_oeb[28] = net80;
 assign io_oeb[2] = net56;
 assign io_oeb[3] = net57;
 assign io_oeb[4] = net58;
 assign io_oeb[5] = net59;
 assign io_oeb[6] = net60;
 assign io_oeb[7] = net61;
 assign io_oeb[8] = net81;
 assign io_oeb[9] = net82;
 assign io_out[10] = net32;
 assign io_out[11] = net33;
 assign io_out[12] = net34;
 assign io_out[13] = net35;
 assign io_out[14] = net36;
 assign io_out[15] = net37;
 assign io_out[16] = net38;
 assign io_out[17] = net39;
 assign io_out[18] = net40;
 assign io_out[19] = net41;
 assign io_out[20] = net42;
 assign io_out[21] = net43;
 assign io_out[22] = net44;
 assign io_out[23] = net45;
 assign io_out[24] = net46;
 assign io_out[25] = net47;
 assign io_out[26] = net48;
 assign io_out[27] = net49;
 assign io_out[28] = net50;
 assign io_out[8] = net30;
 assign io_out[9] = net31;
 assign irq[0] = net51;
 assign irq[1] = net52;
 assign irq[2] = net53;
endmodule

