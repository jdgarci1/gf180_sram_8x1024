magic
tech gf180mcuD
magscale 1 10
timestamp 1702315622
<< obsm1 >>
rect 1344 3076 204736 157442
<< metal2 >>
rect 3808 159264 3920 160064
rect 11424 159264 11536 160064
rect 19040 159264 19152 160064
rect 26656 159264 26768 160064
rect 34272 159264 34384 160064
rect 41888 159264 42000 160064
rect 49504 159264 49616 160064
rect 57120 159264 57232 160064
rect 64736 159264 64848 160064
rect 72352 159264 72464 160064
rect 79968 159264 80080 160064
rect 87584 159264 87696 160064
rect 95200 159264 95312 160064
rect 102816 159264 102928 160064
rect 110432 159264 110544 160064
rect 118048 159264 118160 160064
rect 125664 159264 125776 160064
rect 133280 159264 133392 160064
rect 140896 159264 141008 160064
rect 148512 159264 148624 160064
rect 156128 159264 156240 160064
rect 163744 159264 163856 160064
rect 171360 159264 171472 160064
rect 178976 159264 179088 160064
rect 186592 159264 186704 160064
rect 194208 159264 194320 160064
rect 201824 159264 201936 160064
rect 34272 0 34384 800
rect 102816 0 102928 800
rect 171360 0 171472 800
<< obsm2 >>
rect 1708 159204 3748 159264
rect 3980 159204 11364 159264
rect 11596 159204 18980 159264
rect 19212 159204 26596 159264
rect 26828 159204 34212 159264
rect 34444 159204 41828 159264
rect 42060 159204 49444 159264
rect 49676 159204 57060 159264
rect 57292 159204 64676 159264
rect 64908 159204 72292 159264
rect 72524 159204 79908 159264
rect 80140 159204 87524 159264
rect 87756 159204 95140 159264
rect 95372 159204 102756 159264
rect 102988 159204 110372 159264
rect 110604 159204 117988 159264
rect 118220 159204 125604 159264
rect 125836 159204 133220 159264
rect 133452 159204 140836 159264
rect 141068 159204 148452 159264
rect 148684 159204 156068 159264
rect 156300 159204 163684 159264
rect 163916 159204 171300 159264
rect 171532 159204 178916 159264
rect 179148 159204 186532 159264
rect 186764 159204 194148 159264
rect 194380 159204 201764 159264
rect 201996 159204 204372 159264
rect 1708 860 204372 159204
rect 1708 800 34212 860
rect 34444 800 102756 860
rect 102988 800 171300 860
rect 171532 800 204372 860
<< metal3 >>
rect 0 157920 800 158032
rect 0 154112 800 154224
rect 205332 154112 206132 154224
rect 0 150304 800 150416
rect 0 146496 800 146608
rect 205332 145376 206132 145488
rect 0 142688 800 142800
rect 0 138880 800 138992
rect 205332 136640 206132 136752
rect 0 135072 800 135184
rect 0 131264 800 131376
rect 205332 127904 206132 128016
rect 0 127456 800 127568
rect 0 123648 800 123760
rect 0 119840 800 119952
rect 205332 119168 206132 119280
rect 0 116032 800 116144
rect 0 112224 800 112336
rect 205332 110432 206132 110544
rect 0 108416 800 108528
rect 0 104608 800 104720
rect 205332 101696 206132 101808
rect 0 100800 800 100912
rect 0 96992 800 97104
rect 0 93184 800 93296
rect 205332 92960 206132 93072
rect 0 89376 800 89488
rect 0 85568 800 85680
rect 205332 84224 206132 84336
rect 0 81760 800 81872
rect 0 77952 800 78064
rect 205332 75488 206132 75600
rect 0 74144 800 74256
rect 0 70336 800 70448
rect 205332 66752 206132 66864
rect 0 66528 800 66640
rect 0 62720 800 62832
rect 0 58912 800 59024
rect 205332 58016 206132 58128
rect 0 55104 800 55216
rect 0 51296 800 51408
rect 205332 49280 206132 49392
rect 0 47488 800 47600
rect 0 43680 800 43792
rect 205332 40544 206132 40656
rect 0 39872 800 39984
rect 0 36064 800 36176
rect 0 32256 800 32368
rect 205332 31808 206132 31920
rect 0 28448 800 28560
rect 0 24640 800 24752
rect 205332 23072 206132 23184
rect 0 20832 800 20944
rect 0 17024 800 17136
rect 205332 14336 206132 14448
rect 0 13216 800 13328
rect 0 9408 800 9520
rect 0 5600 800 5712
rect 205332 5600 206132 5712
rect 0 1792 800 1904
<< obsm3 >>
rect 860 157860 205332 158004
rect 800 154284 205332 157860
rect 860 154052 205272 154284
rect 800 150476 205332 154052
rect 860 150244 205332 150476
rect 800 146668 205332 150244
rect 860 146436 205332 146668
rect 800 145548 205332 146436
rect 800 145316 205272 145548
rect 800 142860 205332 145316
rect 860 142628 205332 142860
rect 800 139052 205332 142628
rect 860 138820 205332 139052
rect 800 136812 205332 138820
rect 800 136580 205272 136812
rect 800 135244 205332 136580
rect 860 135012 205332 135244
rect 800 131436 205332 135012
rect 860 131204 205332 131436
rect 800 128076 205332 131204
rect 800 127844 205272 128076
rect 800 127628 205332 127844
rect 860 127396 205332 127628
rect 800 123820 205332 127396
rect 860 123588 205332 123820
rect 800 120012 205332 123588
rect 860 119780 205332 120012
rect 800 119340 205332 119780
rect 800 119108 205272 119340
rect 800 116204 205332 119108
rect 860 115972 205332 116204
rect 800 112396 205332 115972
rect 860 112164 205332 112396
rect 800 110604 205332 112164
rect 800 110372 205272 110604
rect 800 108588 205332 110372
rect 860 108356 205332 108588
rect 800 104780 205332 108356
rect 860 104548 205332 104780
rect 800 101868 205332 104548
rect 800 101636 205272 101868
rect 800 100972 205332 101636
rect 860 100740 205332 100972
rect 800 97164 205332 100740
rect 860 96932 205332 97164
rect 800 93356 205332 96932
rect 860 93132 205332 93356
rect 860 93124 205272 93132
rect 800 92900 205272 93124
rect 800 89548 205332 92900
rect 860 89316 205332 89548
rect 800 85740 205332 89316
rect 860 85508 205332 85740
rect 800 84396 205332 85508
rect 800 84164 205272 84396
rect 800 81932 205332 84164
rect 860 81700 205332 81932
rect 800 78124 205332 81700
rect 860 77892 205332 78124
rect 800 75660 205332 77892
rect 800 75428 205272 75660
rect 800 74316 205332 75428
rect 860 74084 205332 74316
rect 800 70508 205332 74084
rect 860 70276 205332 70508
rect 800 66924 205332 70276
rect 800 66700 205272 66924
rect 860 66692 205272 66700
rect 860 66468 205332 66692
rect 800 62892 205332 66468
rect 860 62660 205332 62892
rect 800 59084 205332 62660
rect 860 58852 205332 59084
rect 800 58188 205332 58852
rect 800 57956 205272 58188
rect 800 55276 205332 57956
rect 860 55044 205332 55276
rect 800 51468 205332 55044
rect 860 51236 205332 51468
rect 800 49452 205332 51236
rect 800 49220 205272 49452
rect 800 47660 205332 49220
rect 860 47428 205332 47660
rect 800 43852 205332 47428
rect 860 43620 205332 43852
rect 800 40716 205332 43620
rect 800 40484 205272 40716
rect 800 40044 205332 40484
rect 860 39812 205332 40044
rect 800 36236 205332 39812
rect 860 36004 205332 36236
rect 800 32428 205332 36004
rect 860 32196 205332 32428
rect 800 31980 205332 32196
rect 800 31748 205272 31980
rect 800 28620 205332 31748
rect 860 28388 205332 28620
rect 800 24812 205332 28388
rect 860 24580 205332 24812
rect 800 23244 205332 24580
rect 800 23012 205272 23244
rect 800 21004 205332 23012
rect 860 20772 205332 21004
rect 800 17196 205332 20772
rect 860 16964 205332 17196
rect 800 14508 205332 16964
rect 800 14276 205272 14508
rect 800 13388 205332 14276
rect 860 13156 205332 13388
rect 800 9580 205332 13156
rect 860 9348 205332 9580
rect 800 5772 205332 9348
rect 860 5540 205272 5772
rect 800 1964 205332 5540
rect 860 1820 205332 1964
<< metal4 >>
rect 4448 3076 4768 156860
rect 5108 3076 5428 156860
rect 35168 3076 35488 156860
rect 35828 3076 36148 156860
rect 65888 142475 66208 156860
rect 66548 34904 66868 156860
rect 96608 39348 96928 156860
rect 97268 34904 97588 156860
rect 127328 34904 127648 156860
rect 65888 3076 66208 20065
rect 66548 3076 66868 20065
rect 96608 3076 96928 17888
rect 97268 3076 97588 21056
rect 127328 3076 127648 21188
rect 127988 3076 128308 156860
rect 158048 3076 158368 156860
rect 158708 3076 159028 156860
rect 188768 3076 189088 156860
rect 189428 3076 189748 156860
<< obsm4 >>
rect 20000 16818 35108 155662
rect 35548 16818 35768 155662
rect 36208 142415 65828 155662
rect 66268 142415 66488 155662
rect 36208 34844 66488 142415
rect 66928 39288 96548 155662
rect 96988 39288 97208 155662
rect 66928 34844 97208 39288
rect 97648 34844 127268 155662
rect 127708 34844 127928 155662
rect 36208 21248 127928 34844
rect 36208 21116 127268 21248
rect 36208 20125 97208 21116
rect 36208 16818 65828 20125
rect 66268 16818 66488 20125
rect 66928 17948 97208 20125
rect 66928 16818 96548 17948
rect 96988 16818 97208 17948
rect 97648 16818 127268 21116
rect 127708 16818 127928 21248
rect 128368 16818 157988 155662
rect 158428 16818 158648 155662
rect 159088 16818 186264 155662
<< metal5 >>
rect 1284 129510 204796 129830
rect 1284 128850 204796 129170
rect 1284 98874 204796 99194
rect 1284 98214 204796 98534
rect 1284 68238 204796 68558
rect 1284 67578 204796 67898
rect 1284 37602 204796 37922
rect 1284 36942 204796 37262
rect 1284 6966 204796 7286
rect 1284 6306 204796 6626
<< labels >>
rlabel metal3 s 205332 5600 206132 5712 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 110432 159264 110544 160064 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 87584 159264 87696 160064 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 64736 159264 64848 160064 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 41888 159264 42000 160064 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 19040 159264 19152 160064 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 157920 800 158032 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 146496 800 146608 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 135072 800 135184 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 123648 800 123760 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 112224 800 112336 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 205332 31808 206132 31920 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 100800 800 100912 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 89376 800 89488 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 77952 800 78064 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 66528 800 66640 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 55104 800 55216 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 43680 800 43792 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 32256 800 32368 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 20832 800 20944 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 9408 800 9520 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 205332 58016 206132 58128 6 io_in[2]
port 22 nsew signal input
rlabel metal3 s 205332 84224 206132 84336 6 io_in[3]
port 23 nsew signal input
rlabel metal3 s 205332 110432 206132 110544 6 io_in[4]
port 24 nsew signal input
rlabel metal3 s 205332 136640 206132 136752 6 io_in[5]
port 25 nsew signal input
rlabel metal2 s 201824 159264 201936 160064 6 io_in[6]
port 26 nsew signal input
rlabel metal2 s 178976 159264 179088 160064 6 io_in[7]
port 27 nsew signal input
rlabel metal2 s 156128 159264 156240 160064 6 io_in[8]
port 28 nsew signal input
rlabel metal2 s 133280 159264 133392 160064 6 io_in[9]
port 29 nsew signal input
rlabel metal3 s 205332 23072 206132 23184 6 io_oeb[0]
port 30 nsew signal output
rlabel metal2 s 95200 159264 95312 160064 6 io_oeb[10]
port 31 nsew signal output
rlabel metal2 s 72352 159264 72464 160064 6 io_oeb[11]
port 32 nsew signal output
rlabel metal2 s 49504 159264 49616 160064 6 io_oeb[12]
port 33 nsew signal output
rlabel metal2 s 26656 159264 26768 160064 6 io_oeb[13]
port 34 nsew signal output
rlabel metal2 s 3808 159264 3920 160064 6 io_oeb[14]
port 35 nsew signal output
rlabel metal3 s 0 150304 800 150416 6 io_oeb[15]
port 36 nsew signal output
rlabel metal3 s 0 138880 800 138992 6 io_oeb[16]
port 37 nsew signal output
rlabel metal3 s 0 127456 800 127568 6 io_oeb[17]
port 38 nsew signal output
rlabel metal3 s 0 116032 800 116144 6 io_oeb[18]
port 39 nsew signal output
rlabel metal3 s 0 104608 800 104720 6 io_oeb[19]
port 40 nsew signal output
rlabel metal3 s 205332 49280 206132 49392 6 io_oeb[1]
port 41 nsew signal output
rlabel metal3 s 0 93184 800 93296 6 io_oeb[20]
port 42 nsew signal output
rlabel metal3 s 0 81760 800 81872 6 io_oeb[21]
port 43 nsew signal output
rlabel metal3 s 0 70336 800 70448 6 io_oeb[22]
port 44 nsew signal output
rlabel metal3 s 0 58912 800 59024 6 io_oeb[23]
port 45 nsew signal output
rlabel metal3 s 0 47488 800 47600 6 io_oeb[24]
port 46 nsew signal output
rlabel metal3 s 0 36064 800 36176 6 io_oeb[25]
port 47 nsew signal output
rlabel metal3 s 0 24640 800 24752 6 io_oeb[26]
port 48 nsew signal output
rlabel metal3 s 0 13216 800 13328 6 io_oeb[27]
port 49 nsew signal output
rlabel metal3 s 0 1792 800 1904 6 io_oeb[28]
port 50 nsew signal output
rlabel metal3 s 205332 75488 206132 75600 6 io_oeb[2]
port 51 nsew signal output
rlabel metal3 s 205332 101696 206132 101808 6 io_oeb[3]
port 52 nsew signal output
rlabel metal3 s 205332 127904 206132 128016 6 io_oeb[4]
port 53 nsew signal output
rlabel metal3 s 205332 154112 206132 154224 6 io_oeb[5]
port 54 nsew signal output
rlabel metal2 s 186592 159264 186704 160064 6 io_oeb[6]
port 55 nsew signal output
rlabel metal2 s 163744 159264 163856 160064 6 io_oeb[7]
port 56 nsew signal output
rlabel metal2 s 140896 159264 141008 160064 6 io_oeb[8]
port 57 nsew signal output
rlabel metal2 s 118048 159264 118160 160064 6 io_oeb[9]
port 58 nsew signal output
rlabel metal3 s 205332 14336 206132 14448 6 io_out[0]
port 59 nsew signal output
rlabel metal2 s 102816 159264 102928 160064 6 io_out[10]
port 60 nsew signal output
rlabel metal2 s 79968 159264 80080 160064 6 io_out[11]
port 61 nsew signal output
rlabel metal2 s 57120 159264 57232 160064 6 io_out[12]
port 62 nsew signal output
rlabel metal2 s 34272 159264 34384 160064 6 io_out[13]
port 63 nsew signal output
rlabel metal2 s 11424 159264 11536 160064 6 io_out[14]
port 64 nsew signal output
rlabel metal3 s 0 154112 800 154224 6 io_out[15]
port 65 nsew signal output
rlabel metal3 s 0 142688 800 142800 6 io_out[16]
port 66 nsew signal output
rlabel metal3 s 0 131264 800 131376 6 io_out[17]
port 67 nsew signal output
rlabel metal3 s 0 119840 800 119952 6 io_out[18]
port 68 nsew signal output
rlabel metal3 s 0 108416 800 108528 6 io_out[19]
port 69 nsew signal output
rlabel metal3 s 205332 40544 206132 40656 6 io_out[1]
port 70 nsew signal output
rlabel metal3 s 0 96992 800 97104 6 io_out[20]
port 71 nsew signal output
rlabel metal3 s 0 85568 800 85680 6 io_out[21]
port 72 nsew signal output
rlabel metal3 s 0 74144 800 74256 6 io_out[22]
port 73 nsew signal output
rlabel metal3 s 0 62720 800 62832 6 io_out[23]
port 74 nsew signal output
rlabel metal3 s 0 51296 800 51408 6 io_out[24]
port 75 nsew signal output
rlabel metal3 s 0 39872 800 39984 6 io_out[25]
port 76 nsew signal output
rlabel metal3 s 0 28448 800 28560 6 io_out[26]
port 77 nsew signal output
rlabel metal3 s 0 17024 800 17136 6 io_out[27]
port 78 nsew signal output
rlabel metal3 s 0 5600 800 5712 6 io_out[28]
port 79 nsew signal output
rlabel metal3 s 205332 66752 206132 66864 6 io_out[2]
port 80 nsew signal output
rlabel metal3 s 205332 92960 206132 93072 6 io_out[3]
port 81 nsew signal output
rlabel metal3 s 205332 119168 206132 119280 6 io_out[4]
port 82 nsew signal output
rlabel metal3 s 205332 145376 206132 145488 6 io_out[5]
port 83 nsew signal output
rlabel metal2 s 194208 159264 194320 160064 6 io_out[6]
port 84 nsew signal output
rlabel metal2 s 171360 159264 171472 160064 6 io_out[7]
port 85 nsew signal output
rlabel metal2 s 148512 159264 148624 160064 6 io_out[8]
port 86 nsew signal output
rlabel metal2 s 125664 159264 125776 160064 6 io_out[9]
port 87 nsew signal output
rlabel metal2 s 34272 0 34384 800 6 irq[0]
port 88 nsew signal output
rlabel metal2 s 102816 0 102928 800 6 irq[1]
port 89 nsew signal output
rlabel metal2 s 171360 0 171472 800 6 irq[2]
port 90 nsew signal output
rlabel metal4 s 4448 3076 4768 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 20065 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 65888 142475 66208 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 17888 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 96608 39348 96928 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 21188 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 127328 34904 127648 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 156860 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 6306 204796 6626 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 36942 204796 37262 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 67578 204796 67898 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 98214 204796 98534 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 128850 204796 129170 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 5108 3076 5428 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 35828 3076 36148 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 66548 3076 66868 20065 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 66548 34904 66868 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 97268 3076 97588 21056 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 97268 34904 97588 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 127988 3076 128308 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 158708 3076 159028 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 189428 3076 189748 156860 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 6966 204796 7286 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 37602 204796 37922 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 68238 204796 68558 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 98874 204796 99194 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 129510 204796 129830 6 vss
port 92 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 206132 160064
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6435020
string GDS_FILE /home/diego/Cinvestav/gf180_sram_8x1024/openlane/user_proj_example/runs/23_12_11_11_24/results/signoff/user_proj_example.magic.gds
string GDS_START 5214300
<< end >>

