magic
tech gf180mcuD
magscale 1 10
timestamp 1702353431
<< obsm1 >>
rect 1344 3076 204848 159570
<< metal2 >>
rect 4032 161772 4144 162572
rect 11648 161772 11760 162572
rect 19264 161772 19376 162572
rect 26880 161772 26992 162572
rect 34496 161772 34608 162572
rect 42112 161772 42224 162572
rect 49728 161772 49840 162572
rect 57344 161772 57456 162572
rect 64960 161772 65072 162572
rect 72576 161772 72688 162572
rect 80192 161772 80304 162572
rect 87808 161772 87920 162572
rect 95424 161772 95536 162572
rect 103040 161772 103152 162572
rect 110656 161772 110768 162572
rect 118272 161772 118384 162572
rect 125888 161772 126000 162572
rect 133504 161772 133616 162572
rect 141120 161772 141232 162572
rect 148736 161772 148848 162572
rect 156352 161772 156464 162572
rect 163968 161772 164080 162572
rect 171584 161772 171696 162572
rect 179200 161772 179312 162572
rect 186816 161772 186928 162572
rect 194432 161772 194544 162572
rect 202048 161772 202160 162572
rect 34272 0 34384 800
rect 103040 0 103152 800
rect 171808 0 171920 800
<< obsm2 >>
rect 1708 161712 3972 161772
rect 4204 161712 11588 161772
rect 11820 161712 19204 161772
rect 19436 161712 26820 161772
rect 27052 161712 34436 161772
rect 34668 161712 42052 161772
rect 42284 161712 49668 161772
rect 49900 161712 57284 161772
rect 57516 161712 64900 161772
rect 65132 161712 72516 161772
rect 72748 161712 80132 161772
rect 80364 161712 87748 161772
rect 87980 161712 95364 161772
rect 95596 161712 102980 161772
rect 103212 161712 110596 161772
rect 110828 161712 118212 161772
rect 118444 161712 125828 161772
rect 126060 161712 133444 161772
rect 133676 161712 141060 161772
rect 141292 161712 148676 161772
rect 148908 161712 156292 161772
rect 156524 161712 163908 161772
rect 164140 161712 171524 161772
rect 171756 161712 179140 161772
rect 179372 161712 186756 161772
rect 186988 161712 194372 161772
rect 194604 161712 201988 161772
rect 202220 161712 204484 161772
rect 1708 860 204484 161712
rect 1708 800 34212 860
rect 34444 800 102980 860
rect 103212 800 171748 860
rect 171980 800 204484 860
<< metal3 >>
rect 0 159264 800 159376
rect 205464 157248 206264 157360
rect 0 155456 800 155568
rect 0 151648 800 151760
rect 205464 148288 206264 148400
rect 0 147840 800 147952
rect 0 144032 800 144144
rect 0 140224 800 140336
rect 205464 139328 206264 139440
rect 0 136416 800 136528
rect 0 132608 800 132720
rect 205464 130368 206264 130480
rect 0 128800 800 128912
rect 0 124992 800 125104
rect 205464 121408 206264 121520
rect 0 121184 800 121296
rect 0 117376 800 117488
rect 0 113568 800 113680
rect 205464 112448 206264 112560
rect 0 109760 800 109872
rect 0 105952 800 106064
rect 205464 103488 206264 103600
rect 0 102144 800 102256
rect 0 98336 800 98448
rect 0 94528 800 94640
rect 205464 94528 206264 94640
rect 0 90720 800 90832
rect 0 86912 800 87024
rect 205464 85568 206264 85680
rect 0 83104 800 83216
rect 0 79296 800 79408
rect 205464 76608 206264 76720
rect 0 75488 800 75600
rect 0 71680 800 71792
rect 0 67872 800 67984
rect 205464 67648 206264 67760
rect 0 64064 800 64176
rect 0 60256 800 60368
rect 205464 58688 206264 58800
rect 0 56448 800 56560
rect 0 52640 800 52752
rect 205464 49728 206264 49840
rect 0 48832 800 48944
rect 0 45024 800 45136
rect 0 41216 800 41328
rect 205464 40768 206264 40880
rect 0 37408 800 37520
rect 0 33600 800 33712
rect 205464 31808 206264 31920
rect 0 29792 800 29904
rect 0 25984 800 26096
rect 205464 22848 206264 22960
rect 0 22176 800 22288
rect 0 18368 800 18480
rect 0 14560 800 14672
rect 205464 13888 206264 14000
rect 0 10752 800 10864
rect 0 6944 800 7056
rect 205464 4928 206264 5040
rect 0 3136 800 3248
<< obsm3 >>
rect 860 159204 205464 159348
rect 800 157420 205464 159204
rect 800 157188 205404 157420
rect 800 155628 205464 157188
rect 860 155396 205464 155628
rect 800 151820 205464 155396
rect 860 151588 205464 151820
rect 800 148460 205464 151588
rect 800 148228 205404 148460
rect 800 148012 205464 148228
rect 860 147780 205464 148012
rect 800 144204 205464 147780
rect 860 143972 205464 144204
rect 800 140396 205464 143972
rect 860 140164 205464 140396
rect 800 139500 205464 140164
rect 800 139268 205404 139500
rect 800 136588 205464 139268
rect 860 136356 205464 136588
rect 800 132780 205464 136356
rect 860 132548 205464 132780
rect 800 130540 205464 132548
rect 800 130308 205404 130540
rect 800 128972 205464 130308
rect 860 128740 205464 128972
rect 800 125164 205464 128740
rect 860 124932 205464 125164
rect 800 121580 205464 124932
rect 800 121356 205404 121580
rect 860 121348 205404 121356
rect 860 121124 205464 121348
rect 800 117548 205464 121124
rect 860 117316 205464 117548
rect 800 113740 205464 117316
rect 860 113508 205464 113740
rect 800 112620 205464 113508
rect 800 112388 205404 112620
rect 800 109932 205464 112388
rect 860 109700 205464 109932
rect 800 106124 205464 109700
rect 860 105892 205464 106124
rect 800 103660 205464 105892
rect 800 103428 205404 103660
rect 800 102316 205464 103428
rect 860 102084 205464 102316
rect 800 98508 205464 102084
rect 860 98276 205464 98508
rect 800 94700 205464 98276
rect 860 94468 205404 94700
rect 800 90892 205464 94468
rect 860 90660 205464 90892
rect 800 87084 205464 90660
rect 860 86852 205464 87084
rect 800 85740 205464 86852
rect 800 85508 205404 85740
rect 800 83276 205464 85508
rect 860 83044 205464 83276
rect 800 79468 205464 83044
rect 860 79236 205464 79468
rect 800 76780 205464 79236
rect 800 76548 205404 76780
rect 800 75660 205464 76548
rect 860 75428 205464 75660
rect 800 71852 205464 75428
rect 860 71620 205464 71852
rect 800 68044 205464 71620
rect 860 67820 205464 68044
rect 860 67812 205404 67820
rect 800 67588 205404 67812
rect 800 64236 205464 67588
rect 860 64004 205464 64236
rect 800 60428 205464 64004
rect 860 60196 205464 60428
rect 800 58860 205464 60196
rect 800 58628 205404 58860
rect 800 56620 205464 58628
rect 860 56388 205464 56620
rect 800 52812 205464 56388
rect 860 52580 205464 52812
rect 800 49900 205464 52580
rect 800 49668 205404 49900
rect 800 49004 205464 49668
rect 860 48772 205464 49004
rect 800 45196 205464 48772
rect 860 44964 205464 45196
rect 800 41388 205464 44964
rect 860 41156 205464 41388
rect 800 40940 205464 41156
rect 800 40708 205404 40940
rect 800 37580 205464 40708
rect 860 37348 205464 37580
rect 800 33772 205464 37348
rect 860 33540 205464 33772
rect 800 31980 205464 33540
rect 800 31748 205404 31980
rect 800 29964 205464 31748
rect 860 29732 205464 29964
rect 800 26156 205464 29732
rect 860 25924 205464 26156
rect 800 23020 205464 25924
rect 800 22788 205404 23020
rect 800 22348 205464 22788
rect 860 22116 205464 22348
rect 800 18540 205464 22116
rect 860 18308 205464 18540
rect 800 14732 205464 18308
rect 860 14500 205464 14732
rect 800 14060 205464 14500
rect 800 13828 205404 14060
rect 800 10924 205464 13828
rect 860 10692 205464 10924
rect 800 7116 205464 10692
rect 860 6884 205464 7116
rect 800 5100 205464 6884
rect 800 4868 205404 5100
rect 800 3308 205464 4868
rect 860 3108 205464 3308
<< metal4 >>
rect 4448 3076 4768 159212
rect 5108 3076 5428 159212
rect 35168 3076 35488 159212
rect 35828 3076 36148 159212
rect 65888 142955 66208 159212
rect 66548 35384 66868 159212
rect 96608 39876 96928 159212
rect 97268 35384 97588 159212
rect 127328 35384 127648 159212
rect 65888 3076 66208 20065
rect 66548 3076 66868 20065
rect 96608 3076 96928 17888
rect 97268 3076 97588 21056
rect 127328 3076 127648 21188
rect 127988 3076 128308 159212
rect 158048 3076 158368 159212
rect 158708 3076 159028 159212
rect 188768 3076 189088 159212
rect 189428 3076 189748 159212
<< obsm4 >>
rect 20000 16818 35108 142572
rect 35548 16818 35768 142572
rect 36208 35324 66488 142572
rect 66928 39816 96548 142572
rect 96988 39816 97208 142572
rect 66928 35324 97208 39816
rect 97648 35324 127268 142572
rect 127708 35324 127928 142572
rect 36208 21248 127928 35324
rect 36208 21116 127268 21248
rect 36208 20125 97208 21116
rect 36208 16818 65828 20125
rect 66268 16818 66488 20125
rect 66928 17948 97208 20125
rect 66928 16818 96548 17948
rect 96988 16818 97208 17948
rect 97648 16818 127268 21116
rect 127708 16818 127928 21248
rect 128368 16818 157988 142572
rect 158428 16818 158648 142572
rect 159088 16818 186264 142572
<< metal5 >>
rect 1284 129510 204908 129830
rect 1284 128850 204908 129170
rect 1284 98874 204908 99194
rect 1284 98214 204908 98534
rect 1284 68238 204908 68558
rect 1284 67578 204908 67898
rect 1284 37602 204908 37922
rect 1284 36942 204908 37262
rect 1284 6966 204908 7286
rect 1284 6306 204908 6626
<< labels >>
rlabel metal3 s 205464 4928 206264 5040 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 110656 161772 110768 162572 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 87808 161772 87920 162572 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 64960 161772 65072 162572 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 42112 161772 42224 162572 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 19264 161772 19376 162572 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 159264 800 159376 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 147840 800 147952 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 136416 800 136528 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 124992 800 125104 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 113568 800 113680 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 205464 31808 206264 31920 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 102144 800 102256 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 90720 800 90832 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 79296 800 79408 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 67872 800 67984 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 56448 800 56560 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 45024 800 45136 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 33600 800 33712 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 22176 800 22288 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 10752 800 10864 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 205464 58688 206264 58800 6 io_in[2]
port 22 nsew signal input
rlabel metal3 s 205464 85568 206264 85680 6 io_in[3]
port 23 nsew signal input
rlabel metal3 s 205464 112448 206264 112560 6 io_in[4]
port 24 nsew signal input
rlabel metal3 s 205464 139328 206264 139440 6 io_in[5]
port 25 nsew signal input
rlabel metal2 s 202048 161772 202160 162572 6 io_in[6]
port 26 nsew signal input
rlabel metal2 s 179200 161772 179312 162572 6 io_in[7]
port 27 nsew signal input
rlabel metal2 s 156352 161772 156464 162572 6 io_in[8]
port 28 nsew signal input
rlabel metal2 s 133504 161772 133616 162572 6 io_in[9]
port 29 nsew signal input
rlabel metal3 s 205464 22848 206264 22960 6 io_oeb[0]
port 30 nsew signal output
rlabel metal2 s 95424 161772 95536 162572 6 io_oeb[10]
port 31 nsew signal output
rlabel metal2 s 72576 161772 72688 162572 6 io_oeb[11]
port 32 nsew signal output
rlabel metal2 s 49728 161772 49840 162572 6 io_oeb[12]
port 33 nsew signal output
rlabel metal2 s 26880 161772 26992 162572 6 io_oeb[13]
port 34 nsew signal output
rlabel metal2 s 4032 161772 4144 162572 6 io_oeb[14]
port 35 nsew signal output
rlabel metal3 s 0 151648 800 151760 6 io_oeb[15]
port 36 nsew signal output
rlabel metal3 s 0 140224 800 140336 6 io_oeb[16]
port 37 nsew signal output
rlabel metal3 s 0 128800 800 128912 6 io_oeb[17]
port 38 nsew signal output
rlabel metal3 s 0 117376 800 117488 6 io_oeb[18]
port 39 nsew signal output
rlabel metal3 s 0 105952 800 106064 6 io_oeb[19]
port 40 nsew signal output
rlabel metal3 s 205464 49728 206264 49840 6 io_oeb[1]
port 41 nsew signal output
rlabel metal3 s 0 94528 800 94640 6 io_oeb[20]
port 42 nsew signal output
rlabel metal3 s 0 83104 800 83216 6 io_oeb[21]
port 43 nsew signal output
rlabel metal3 s 0 71680 800 71792 6 io_oeb[22]
port 44 nsew signal output
rlabel metal3 s 0 60256 800 60368 6 io_oeb[23]
port 45 nsew signal output
rlabel metal3 s 0 48832 800 48944 6 io_oeb[24]
port 46 nsew signal output
rlabel metal3 s 0 37408 800 37520 6 io_oeb[25]
port 47 nsew signal output
rlabel metal3 s 0 25984 800 26096 6 io_oeb[26]
port 48 nsew signal output
rlabel metal3 s 0 14560 800 14672 6 io_oeb[27]
port 49 nsew signal output
rlabel metal3 s 0 3136 800 3248 6 io_oeb[28]
port 50 nsew signal output
rlabel metal3 s 205464 76608 206264 76720 6 io_oeb[2]
port 51 nsew signal output
rlabel metal3 s 205464 103488 206264 103600 6 io_oeb[3]
port 52 nsew signal output
rlabel metal3 s 205464 130368 206264 130480 6 io_oeb[4]
port 53 nsew signal output
rlabel metal3 s 205464 157248 206264 157360 6 io_oeb[5]
port 54 nsew signal output
rlabel metal2 s 186816 161772 186928 162572 6 io_oeb[6]
port 55 nsew signal output
rlabel metal2 s 163968 161772 164080 162572 6 io_oeb[7]
port 56 nsew signal output
rlabel metal2 s 141120 161772 141232 162572 6 io_oeb[8]
port 57 nsew signal output
rlabel metal2 s 118272 161772 118384 162572 6 io_oeb[9]
port 58 nsew signal output
rlabel metal3 s 205464 13888 206264 14000 6 io_out[0]
port 59 nsew signal output
rlabel metal2 s 103040 161772 103152 162572 6 io_out[10]
port 60 nsew signal output
rlabel metal2 s 80192 161772 80304 162572 6 io_out[11]
port 61 nsew signal output
rlabel metal2 s 57344 161772 57456 162572 6 io_out[12]
port 62 nsew signal output
rlabel metal2 s 34496 161772 34608 162572 6 io_out[13]
port 63 nsew signal output
rlabel metal2 s 11648 161772 11760 162572 6 io_out[14]
port 64 nsew signal output
rlabel metal3 s 0 155456 800 155568 6 io_out[15]
port 65 nsew signal output
rlabel metal3 s 0 144032 800 144144 6 io_out[16]
port 66 nsew signal output
rlabel metal3 s 0 132608 800 132720 6 io_out[17]
port 67 nsew signal output
rlabel metal3 s 0 121184 800 121296 6 io_out[18]
port 68 nsew signal output
rlabel metal3 s 0 109760 800 109872 6 io_out[19]
port 69 nsew signal output
rlabel metal3 s 205464 40768 206264 40880 6 io_out[1]
port 70 nsew signal output
rlabel metal3 s 0 98336 800 98448 6 io_out[20]
port 71 nsew signal output
rlabel metal3 s 0 86912 800 87024 6 io_out[21]
port 72 nsew signal output
rlabel metal3 s 0 75488 800 75600 6 io_out[22]
port 73 nsew signal output
rlabel metal3 s 0 64064 800 64176 6 io_out[23]
port 74 nsew signal output
rlabel metal3 s 0 52640 800 52752 6 io_out[24]
port 75 nsew signal output
rlabel metal3 s 0 41216 800 41328 6 io_out[25]
port 76 nsew signal output
rlabel metal3 s 0 29792 800 29904 6 io_out[26]
port 77 nsew signal output
rlabel metal3 s 0 18368 800 18480 6 io_out[27]
port 78 nsew signal output
rlabel metal3 s 0 6944 800 7056 6 io_out[28]
port 79 nsew signal output
rlabel metal3 s 205464 67648 206264 67760 6 io_out[2]
port 80 nsew signal output
rlabel metal3 s 205464 94528 206264 94640 6 io_out[3]
port 81 nsew signal output
rlabel metal3 s 205464 121408 206264 121520 6 io_out[4]
port 82 nsew signal output
rlabel metal3 s 205464 148288 206264 148400 6 io_out[5]
port 83 nsew signal output
rlabel metal2 s 194432 161772 194544 162572 6 io_out[6]
port 84 nsew signal output
rlabel metal2 s 171584 161772 171696 162572 6 io_out[7]
port 85 nsew signal output
rlabel metal2 s 148736 161772 148848 162572 6 io_out[8]
port 86 nsew signal output
rlabel metal2 s 125888 161772 126000 162572 6 io_out[9]
port 87 nsew signal output
rlabel metal2 s 34272 0 34384 800 6 irq[0]
port 88 nsew signal output
rlabel metal2 s 103040 0 103152 800 6 irq[1]
port 89 nsew signal output
rlabel metal2 s 171808 0 171920 800 6 irq[2]
port 90 nsew signal output
rlabel metal4 s 4448 3076 4768 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 20065 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 65888 142955 66208 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 17888 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 96608 39876 96928 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 21188 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 127328 35384 127648 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 159212 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 6306 204908 6626 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 36942 204908 37262 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 67578 204908 67898 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 98214 204908 98534 6 vdd
port 91 nsew power bidirectional
rlabel metal5 s 1284 128850 204908 129170 6 vdd
port 91 nsew power bidirectional
rlabel metal4 s 5108 3076 5428 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 35828 3076 36148 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 66548 3076 66868 20065 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 66548 35384 66868 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 97268 3076 97588 21056 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 97268 35384 97588 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 127988 3076 128308 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 158708 3076 159028 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal4 s 189428 3076 189748 159212 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 6966 204908 7286 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 37602 204908 37922 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 68238 204908 68558 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 98874 204908 99194 6 vss
port 92 nsew ground bidirectional
rlabel metal5 s 1284 129510 204908 129830 6 vss
port 92 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 206264 162572
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6411298
string GDS_FILE /home/diego/Cinvestav/gf180_sram_8x1024/openlane/user_proj_example/runs/23_12_11_21_53/results/signoff/user_proj_example.magic.gds
string GDS_START 5160914
<< end >>

