VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1031.320 BY 812.860 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 24.640 1031.320 25.200 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 808.860 553.840 812.860 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 808.860 439.600 812.860 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 808.860 325.360 812.860 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 808.860 211.120 812.860 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 808.860 96.880 812.860 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 796.320 4.000 796.880 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.200 4.000 739.760 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 159.040 1031.320 159.600 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 396.480 4.000 397.040 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.360 4.000 339.920 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.240 4.000 282.800 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END io_in[28]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 293.440 1031.320 294.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 427.840 1031.320 428.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 562.240 1031.320 562.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 696.640 1031.320 697.200 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 808.860 1010.800 812.860 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 896.000 808.860 896.560 812.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 808.860 782.320 812.860 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 667.520 808.860 668.080 812.860 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 114.240 1031.320 114.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 808.860 477.680 812.860 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 808.860 363.440 812.860 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 808.860 249.200 812.860 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 808.860 134.960 812.860 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 808.860 20.720 812.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 758.240 4.000 758.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 701.120 4.000 701.680 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 644.000 4.000 644.560 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 586.880 4.000 587.440 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 529.760 4.000 530.320 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 248.640 1031.320 249.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.640 4.000 473.200 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 415.520 4.000 416.080 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.280 4.000 301.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.160 4.000 244.720 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 4.000 187.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 4.000 16.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 383.040 1031.320 383.600 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 517.440 1031.320 518.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 651.840 1031.320 652.400 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 786.240 1031.320 786.800 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 808.860 934.640 812.860 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 808.860 820.400 812.860 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 808.860 706.160 812.860 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 808.860 591.920 812.860 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 69.440 1031.320 70.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 808.860 515.760 812.860 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 808.860 401.520 812.860 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 808.860 287.280 812.860 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 808.860 173.040 812.860 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 808.860 58.800 812.860 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 777.280 4.000 777.840 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 720.160 4.000 720.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.040 4.000 663.600 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 605.920 4.000 606.480 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 203.840 1031.320 204.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.680 4.000 492.240 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 434.560 4.000 435.120 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.440 4.000 378.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 4.000 92.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END io_out[28]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 338.240 1031.320 338.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 472.640 1031.320 473.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 607.040 1031.320 607.600 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1027.320 741.440 1031.320 742.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 972.160 808.860 972.720 812.860 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 808.860 858.480 812.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 808.860 744.240 812.860 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 808.860 630.000 812.860 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 859.040 0.000 859.600 4.000 ;
    END
  END irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 100.325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 714.775 331.040 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 89.440 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 199.380 484.640 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 105.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 176.920 638.240 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 796.060 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 25.540 15.380 27.140 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 15.380 180.740 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 15.380 334.340 100.325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 176.920 334.340 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 15.380 487.940 105.280 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 176.920 487.940 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.940 15.380 641.540 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 793.540 15.380 795.140 796.060 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 947.140 15.380 948.740 796.060 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1024.240 797.850 ;
      LAYER Metal2 ;
        RECT 8.540 808.560 19.860 808.860 ;
        RECT 21.020 808.560 57.940 808.860 ;
        RECT 59.100 808.560 96.020 808.860 ;
        RECT 97.180 808.560 134.100 808.860 ;
        RECT 135.260 808.560 172.180 808.860 ;
        RECT 173.340 808.560 210.260 808.860 ;
        RECT 211.420 808.560 248.340 808.860 ;
        RECT 249.500 808.560 286.420 808.860 ;
        RECT 287.580 808.560 324.500 808.860 ;
        RECT 325.660 808.560 362.580 808.860 ;
        RECT 363.740 808.560 400.660 808.860 ;
        RECT 401.820 808.560 438.740 808.860 ;
        RECT 439.900 808.560 476.820 808.860 ;
        RECT 477.980 808.560 514.900 808.860 ;
        RECT 516.060 808.560 552.980 808.860 ;
        RECT 554.140 808.560 591.060 808.860 ;
        RECT 592.220 808.560 629.140 808.860 ;
        RECT 630.300 808.560 667.220 808.860 ;
        RECT 668.380 808.560 705.300 808.860 ;
        RECT 706.460 808.560 743.380 808.860 ;
        RECT 744.540 808.560 781.460 808.860 ;
        RECT 782.620 808.560 819.540 808.860 ;
        RECT 820.700 808.560 857.620 808.860 ;
        RECT 858.780 808.560 895.700 808.860 ;
        RECT 896.860 808.560 933.780 808.860 ;
        RECT 934.940 808.560 971.860 808.860 ;
        RECT 973.020 808.560 1009.940 808.860 ;
        RECT 1011.100 808.560 1022.420 808.860 ;
        RECT 8.540 4.300 1022.420 808.560 ;
        RECT 8.540 4.000 171.060 4.300 ;
        RECT 172.220 4.000 514.900 4.300 ;
        RECT 516.060 4.000 858.740 4.300 ;
        RECT 859.900 4.000 1022.420 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 796.020 1027.320 796.740 ;
        RECT 4.000 787.100 1027.320 796.020 ;
        RECT 4.000 785.940 1027.020 787.100 ;
        RECT 4.000 778.140 1027.320 785.940 ;
        RECT 4.300 776.980 1027.320 778.140 ;
        RECT 4.000 759.100 1027.320 776.980 ;
        RECT 4.300 757.940 1027.320 759.100 ;
        RECT 4.000 742.300 1027.320 757.940 ;
        RECT 4.000 741.140 1027.020 742.300 ;
        RECT 4.000 740.060 1027.320 741.140 ;
        RECT 4.300 738.900 1027.320 740.060 ;
        RECT 4.000 721.020 1027.320 738.900 ;
        RECT 4.300 719.860 1027.320 721.020 ;
        RECT 4.000 701.980 1027.320 719.860 ;
        RECT 4.300 700.820 1027.320 701.980 ;
        RECT 4.000 697.500 1027.320 700.820 ;
        RECT 4.000 696.340 1027.020 697.500 ;
        RECT 4.000 682.940 1027.320 696.340 ;
        RECT 4.300 681.780 1027.320 682.940 ;
        RECT 4.000 663.900 1027.320 681.780 ;
        RECT 4.300 662.740 1027.320 663.900 ;
        RECT 4.000 652.700 1027.320 662.740 ;
        RECT 4.000 651.540 1027.020 652.700 ;
        RECT 4.000 644.860 1027.320 651.540 ;
        RECT 4.300 643.700 1027.320 644.860 ;
        RECT 4.000 625.820 1027.320 643.700 ;
        RECT 4.300 624.660 1027.320 625.820 ;
        RECT 4.000 607.900 1027.320 624.660 ;
        RECT 4.000 606.780 1027.020 607.900 ;
        RECT 4.300 606.740 1027.020 606.780 ;
        RECT 4.300 605.620 1027.320 606.740 ;
        RECT 4.000 587.740 1027.320 605.620 ;
        RECT 4.300 586.580 1027.320 587.740 ;
        RECT 4.000 568.700 1027.320 586.580 ;
        RECT 4.300 567.540 1027.320 568.700 ;
        RECT 4.000 563.100 1027.320 567.540 ;
        RECT 4.000 561.940 1027.020 563.100 ;
        RECT 4.000 549.660 1027.320 561.940 ;
        RECT 4.300 548.500 1027.320 549.660 ;
        RECT 4.000 530.620 1027.320 548.500 ;
        RECT 4.300 529.460 1027.320 530.620 ;
        RECT 4.000 518.300 1027.320 529.460 ;
        RECT 4.000 517.140 1027.020 518.300 ;
        RECT 4.000 511.580 1027.320 517.140 ;
        RECT 4.300 510.420 1027.320 511.580 ;
        RECT 4.000 492.540 1027.320 510.420 ;
        RECT 4.300 491.380 1027.320 492.540 ;
        RECT 4.000 473.500 1027.320 491.380 ;
        RECT 4.300 472.340 1027.020 473.500 ;
        RECT 4.000 454.460 1027.320 472.340 ;
        RECT 4.300 453.300 1027.320 454.460 ;
        RECT 4.000 435.420 1027.320 453.300 ;
        RECT 4.300 434.260 1027.320 435.420 ;
        RECT 4.000 428.700 1027.320 434.260 ;
        RECT 4.000 427.540 1027.020 428.700 ;
        RECT 4.000 416.380 1027.320 427.540 ;
        RECT 4.300 415.220 1027.320 416.380 ;
        RECT 4.000 397.340 1027.320 415.220 ;
        RECT 4.300 396.180 1027.320 397.340 ;
        RECT 4.000 383.900 1027.320 396.180 ;
        RECT 4.000 382.740 1027.020 383.900 ;
        RECT 4.000 378.300 1027.320 382.740 ;
        RECT 4.300 377.140 1027.320 378.300 ;
        RECT 4.000 359.260 1027.320 377.140 ;
        RECT 4.300 358.100 1027.320 359.260 ;
        RECT 4.000 340.220 1027.320 358.100 ;
        RECT 4.300 339.100 1027.320 340.220 ;
        RECT 4.300 339.060 1027.020 339.100 ;
        RECT 4.000 337.940 1027.020 339.060 ;
        RECT 4.000 321.180 1027.320 337.940 ;
        RECT 4.300 320.020 1027.320 321.180 ;
        RECT 4.000 302.140 1027.320 320.020 ;
        RECT 4.300 300.980 1027.320 302.140 ;
        RECT 4.000 294.300 1027.320 300.980 ;
        RECT 4.000 293.140 1027.020 294.300 ;
        RECT 4.000 283.100 1027.320 293.140 ;
        RECT 4.300 281.940 1027.320 283.100 ;
        RECT 4.000 264.060 1027.320 281.940 ;
        RECT 4.300 262.900 1027.320 264.060 ;
        RECT 4.000 249.500 1027.320 262.900 ;
        RECT 4.000 248.340 1027.020 249.500 ;
        RECT 4.000 245.020 1027.320 248.340 ;
        RECT 4.300 243.860 1027.320 245.020 ;
        RECT 4.000 225.980 1027.320 243.860 ;
        RECT 4.300 224.820 1027.320 225.980 ;
        RECT 4.000 206.940 1027.320 224.820 ;
        RECT 4.300 205.780 1027.320 206.940 ;
        RECT 4.000 204.700 1027.320 205.780 ;
        RECT 4.000 203.540 1027.020 204.700 ;
        RECT 4.000 187.900 1027.320 203.540 ;
        RECT 4.300 186.740 1027.320 187.900 ;
        RECT 4.000 168.860 1027.320 186.740 ;
        RECT 4.300 167.700 1027.320 168.860 ;
        RECT 4.000 159.900 1027.320 167.700 ;
        RECT 4.000 158.740 1027.020 159.900 ;
        RECT 4.000 149.820 1027.320 158.740 ;
        RECT 4.300 148.660 1027.320 149.820 ;
        RECT 4.000 130.780 1027.320 148.660 ;
        RECT 4.300 129.620 1027.320 130.780 ;
        RECT 4.000 115.100 1027.320 129.620 ;
        RECT 4.000 113.940 1027.020 115.100 ;
        RECT 4.000 111.740 1027.320 113.940 ;
        RECT 4.300 110.580 1027.320 111.740 ;
        RECT 4.000 92.700 1027.320 110.580 ;
        RECT 4.300 91.540 1027.320 92.700 ;
        RECT 4.000 73.660 1027.320 91.540 ;
        RECT 4.300 72.500 1027.320 73.660 ;
        RECT 4.000 70.300 1027.320 72.500 ;
        RECT 4.000 69.140 1027.020 70.300 ;
        RECT 4.000 54.620 1027.320 69.140 ;
        RECT 4.300 53.460 1027.320 54.620 ;
        RECT 4.000 35.580 1027.320 53.460 ;
        RECT 4.300 34.420 1027.320 35.580 ;
        RECT 4.000 25.500 1027.320 34.420 ;
        RECT 4.000 24.340 1027.020 25.500 ;
        RECT 4.000 16.540 1027.320 24.340 ;
        RECT 4.300 15.540 1027.320 16.540 ;
      LAYER Metal4 ;
        RECT 100.000 84.090 175.540 712.860 ;
        RECT 177.740 84.090 178.840 712.860 ;
        RECT 181.040 176.620 332.440 712.860 ;
        RECT 334.640 199.080 482.740 712.860 ;
        RECT 484.940 199.080 486.040 712.860 ;
        RECT 334.640 176.620 486.040 199.080 ;
        RECT 488.240 176.620 636.340 712.860 ;
        RECT 638.540 176.620 639.640 712.860 ;
        RECT 181.040 106.240 639.640 176.620 ;
        RECT 181.040 105.580 636.340 106.240 ;
        RECT 181.040 100.625 486.040 105.580 ;
        RECT 181.040 84.090 329.140 100.625 ;
        RECT 331.340 84.090 332.440 100.625 ;
        RECT 334.640 89.740 486.040 100.625 ;
        RECT 334.640 84.090 482.740 89.740 ;
        RECT 484.940 84.090 486.040 89.740 ;
        RECT 488.240 84.090 636.340 105.580 ;
        RECT 638.540 84.090 639.640 106.240 ;
        RECT 641.840 84.090 789.940 712.860 ;
        RECT 792.140 84.090 793.240 712.860 ;
        RECT 795.440 84.090 931.320 712.860 ;
  END
END user_proj_example
END LIBRARY

