magic
tech gf180mcuD
magscale 1 10
timestamp 1702321784
<< metal1 >>
rect 133298 157390 133310 157442
rect 133362 157439 133374 157442
rect 134194 157439 134206 157442
rect 133362 157393 134206 157439
rect 133362 157390 133374 157393
rect 134194 157390 134206 157393
rect 134258 157390 134270 157442
rect 87602 157054 87614 157106
rect 87666 157103 87678 157106
rect 88498 157103 88510 157106
rect 87666 157057 88510 157103
rect 87666 157054 87678 157057
rect 88498 157054 88510 157057
rect 88562 157103 88574 157106
rect 89394 157103 89406 157106
rect 88562 157057 89406 157103
rect 88562 157054 88574 157057
rect 89394 157054 89406 157057
rect 89458 157054 89470 157106
rect 156258 157054 156270 157106
rect 156322 157103 156334 157106
rect 157042 157103 157054 157106
rect 156322 157057 157054 157103
rect 156322 157054 156334 157057
rect 157042 157054 157054 157057
rect 157106 157103 157118 157106
rect 157938 157103 157950 157106
rect 157106 157057 157950 157103
rect 157106 157054 157118 157057
rect 157938 157054 157950 157057
rect 158002 157054 158014 157106
rect 1344 156826 204736 156860
rect 1344 156774 5138 156826
rect 5190 156774 5242 156826
rect 5294 156774 5346 156826
rect 5398 156774 35858 156826
rect 35910 156774 35962 156826
rect 36014 156774 36066 156826
rect 36118 156774 66578 156826
rect 66630 156774 66682 156826
rect 66734 156774 66786 156826
rect 66838 156774 97298 156826
rect 97350 156774 97402 156826
rect 97454 156774 97506 156826
rect 97558 156774 128018 156826
rect 128070 156774 128122 156826
rect 128174 156774 128226 156826
rect 128278 156774 158738 156826
rect 158790 156774 158842 156826
rect 158894 156774 158946 156826
rect 158998 156774 189458 156826
rect 189510 156774 189562 156826
rect 189614 156774 189666 156826
rect 189718 156774 204736 156826
rect 1344 156740 204736 156774
rect 11678 156658 11730 156670
rect 11678 156594 11730 156606
rect 19070 156658 19122 156670
rect 19070 156594 19122 156606
rect 19294 156658 19346 156670
rect 19294 156594 19346 156606
rect 34526 156658 34578 156670
rect 34526 156594 34578 156606
rect 43710 156658 43762 156670
rect 43710 156594 43762 156606
rect 57374 156658 57426 156670
rect 57374 156594 57426 156606
rect 66558 156658 66610 156670
rect 66558 156594 66610 156606
rect 80222 156658 80274 156670
rect 80222 156594 80274 156606
rect 89406 156658 89458 156670
rect 89406 156594 89458 156606
rect 103070 156658 103122 156670
rect 103070 156594 103122 156606
rect 110462 156658 110514 156670
rect 110462 156594 110514 156606
rect 110686 156658 110738 156670
rect 110686 156594 110738 156606
rect 125918 156658 125970 156670
rect 125918 156594 125970 156606
rect 135102 156658 135154 156670
rect 135102 156594 135154 156606
rect 148766 156658 148818 156670
rect 148766 156594 148818 156606
rect 157950 156658 158002 156670
rect 157950 156594 158002 156606
rect 163998 156658 164050 156670
rect 163998 156594 164050 156606
rect 186846 156658 186898 156670
rect 186846 156594 186898 156606
rect 1698 156494 1710 156546
rect 1762 156494 1774 156546
rect 87602 156494 87614 156546
rect 87666 156494 87678 156546
rect 41906 156382 41918 156434
rect 41970 156382 41982 156434
rect 64754 156382 64766 156434
rect 64818 156382 64830 156434
rect 88498 156382 88510 156434
rect 88562 156382 88574 156434
rect 134194 156382 134206 156434
rect 134258 156382 134270 156434
rect 157042 156382 157054 156434
rect 157106 156382 157118 156434
rect 2370 156270 2382 156322
rect 2434 156270 2446 156322
rect 20066 156270 20078 156322
rect 20130 156270 20142 156322
rect 42802 156270 42814 156322
rect 42866 156270 42878 156322
rect 65314 156270 65326 156322
rect 65378 156270 65390 156322
rect 111122 156270 111134 156322
rect 111186 156270 111198 156322
rect 156370 156270 156382 156322
rect 156434 156270 156446 156322
rect 4062 156210 4114 156222
rect 4062 156146 4114 156158
rect 26910 156210 26962 156222
rect 26910 156146 26962 156158
rect 49758 156210 49810 156222
rect 49758 156146 49810 156158
rect 72606 156210 72658 156222
rect 72606 156146 72658 156158
rect 95454 156210 95506 156222
rect 95454 156146 95506 156158
rect 118302 156210 118354 156222
rect 118302 156146 118354 156158
rect 133422 156210 133474 156222
rect 133422 156146 133474 156158
rect 141150 156210 141202 156222
rect 141150 156146 141202 156158
rect 1344 156042 204736 156076
rect 1344 155990 4478 156042
rect 4530 155990 4582 156042
rect 4634 155990 4686 156042
rect 4738 155990 35198 156042
rect 35250 155990 35302 156042
rect 35354 155990 35406 156042
rect 35458 155990 65918 156042
rect 65970 155990 66022 156042
rect 66074 155990 66126 156042
rect 66178 155990 96638 156042
rect 96690 155990 96742 156042
rect 96794 155990 96846 156042
rect 96898 155990 127358 156042
rect 127410 155990 127462 156042
rect 127514 155990 127566 156042
rect 127618 155990 158078 156042
rect 158130 155990 158182 156042
rect 158234 155990 158286 156042
rect 158338 155990 188798 156042
rect 188850 155990 188902 156042
rect 188954 155990 189006 156042
rect 189058 155990 204736 156042
rect 1344 155956 204736 155990
rect 171838 155874 171890 155886
rect 171838 155810 171890 155822
rect 1822 155762 1874 155774
rect 194898 155710 194910 155762
rect 194962 155710 194974 155762
rect 1822 155698 1874 155710
rect 174178 155598 174190 155650
rect 174242 155598 174254 155650
rect 196578 155598 196590 155650
rect 196642 155598 196654 155650
rect 174638 155426 174690 155438
rect 174638 155362 174690 155374
rect 197486 155426 197538 155438
rect 197486 155362 197538 155374
rect 1344 155258 204736 155292
rect 1344 155206 5138 155258
rect 5190 155206 5242 155258
rect 5294 155206 5346 155258
rect 5398 155206 35858 155258
rect 35910 155206 35962 155258
rect 36014 155206 36066 155258
rect 36118 155206 66578 155258
rect 66630 155206 66682 155258
rect 66734 155206 66786 155258
rect 66838 155206 97298 155258
rect 97350 155206 97402 155258
rect 97454 155206 97506 155258
rect 97558 155206 128018 155258
rect 128070 155206 128122 155258
rect 128174 155206 128226 155258
rect 128278 155206 158738 155258
rect 158790 155206 158842 155258
rect 158894 155206 158946 155258
rect 158998 155206 189458 155258
rect 189510 155206 189562 155258
rect 189614 155206 189666 155258
rect 189718 155206 204736 155258
rect 1344 155172 204736 155206
rect 1710 154978 1762 154990
rect 1710 154914 1762 154926
rect 204318 154978 204370 154990
rect 204318 154914 204370 154926
rect 1344 154474 204736 154508
rect 1344 154422 4478 154474
rect 4530 154422 4582 154474
rect 4634 154422 4686 154474
rect 4738 154422 35198 154474
rect 35250 154422 35302 154474
rect 35354 154422 35406 154474
rect 35458 154422 65918 154474
rect 65970 154422 66022 154474
rect 66074 154422 66126 154474
rect 66178 154422 96638 154474
rect 96690 154422 96742 154474
rect 96794 154422 96846 154474
rect 96898 154422 127358 154474
rect 127410 154422 127462 154474
rect 127514 154422 127566 154474
rect 127618 154422 158078 154474
rect 158130 154422 158182 154474
rect 158234 154422 158286 154474
rect 158338 154422 188798 154474
rect 188850 154422 188902 154474
rect 188954 154422 189006 154474
rect 189058 154422 204736 154474
rect 1344 154388 204736 154422
rect 1344 153690 204736 153724
rect 1344 153638 5138 153690
rect 5190 153638 5242 153690
rect 5294 153638 5346 153690
rect 5398 153638 35858 153690
rect 35910 153638 35962 153690
rect 36014 153638 36066 153690
rect 36118 153638 66578 153690
rect 66630 153638 66682 153690
rect 66734 153638 66786 153690
rect 66838 153638 97298 153690
rect 97350 153638 97402 153690
rect 97454 153638 97506 153690
rect 97558 153638 128018 153690
rect 128070 153638 128122 153690
rect 128174 153638 128226 153690
rect 128278 153638 158738 153690
rect 158790 153638 158842 153690
rect 158894 153638 158946 153690
rect 158998 153638 189458 153690
rect 189510 153638 189562 153690
rect 189614 153638 189666 153690
rect 189718 153638 204736 153690
rect 1344 153604 204736 153638
rect 1344 152906 204736 152940
rect 1344 152854 4478 152906
rect 4530 152854 4582 152906
rect 4634 152854 4686 152906
rect 4738 152854 35198 152906
rect 35250 152854 35302 152906
rect 35354 152854 35406 152906
rect 35458 152854 65918 152906
rect 65970 152854 66022 152906
rect 66074 152854 66126 152906
rect 66178 152854 96638 152906
rect 96690 152854 96742 152906
rect 96794 152854 96846 152906
rect 96898 152854 127358 152906
rect 127410 152854 127462 152906
rect 127514 152854 127566 152906
rect 127618 152854 158078 152906
rect 158130 152854 158182 152906
rect 158234 152854 158286 152906
rect 158338 152854 188798 152906
rect 188850 152854 188902 152906
rect 188954 152854 189006 152906
rect 189058 152854 204736 152906
rect 1344 152820 204736 152854
rect 1344 152122 204736 152156
rect 1344 152070 5138 152122
rect 5190 152070 5242 152122
rect 5294 152070 5346 152122
rect 5398 152070 35858 152122
rect 35910 152070 35962 152122
rect 36014 152070 36066 152122
rect 36118 152070 66578 152122
rect 66630 152070 66682 152122
rect 66734 152070 66786 152122
rect 66838 152070 97298 152122
rect 97350 152070 97402 152122
rect 97454 152070 97506 152122
rect 97558 152070 128018 152122
rect 128070 152070 128122 152122
rect 128174 152070 128226 152122
rect 128278 152070 158738 152122
rect 158790 152070 158842 152122
rect 158894 152070 158946 152122
rect 158998 152070 189458 152122
rect 189510 152070 189562 152122
rect 189614 152070 189666 152122
rect 189718 152070 204736 152122
rect 1344 152036 204736 152070
rect 1344 151338 204736 151372
rect 1344 151286 4478 151338
rect 4530 151286 4582 151338
rect 4634 151286 4686 151338
rect 4738 151286 35198 151338
rect 35250 151286 35302 151338
rect 35354 151286 35406 151338
rect 35458 151286 65918 151338
rect 65970 151286 66022 151338
rect 66074 151286 66126 151338
rect 66178 151286 96638 151338
rect 96690 151286 96742 151338
rect 96794 151286 96846 151338
rect 96898 151286 127358 151338
rect 127410 151286 127462 151338
rect 127514 151286 127566 151338
rect 127618 151286 158078 151338
rect 158130 151286 158182 151338
rect 158234 151286 158286 151338
rect 158338 151286 188798 151338
rect 188850 151286 188902 151338
rect 188954 151286 189006 151338
rect 189058 151286 204736 151338
rect 1344 151252 204736 151286
rect 1710 151058 1762 151070
rect 1710 150994 1762 151006
rect 1344 150554 204736 150588
rect 1344 150502 5138 150554
rect 5190 150502 5242 150554
rect 5294 150502 5346 150554
rect 5398 150502 35858 150554
rect 35910 150502 35962 150554
rect 36014 150502 36066 150554
rect 36118 150502 66578 150554
rect 66630 150502 66682 150554
rect 66734 150502 66786 150554
rect 66838 150502 97298 150554
rect 97350 150502 97402 150554
rect 97454 150502 97506 150554
rect 97558 150502 128018 150554
rect 128070 150502 128122 150554
rect 128174 150502 128226 150554
rect 128278 150502 158738 150554
rect 158790 150502 158842 150554
rect 158894 150502 158946 150554
rect 158998 150502 189458 150554
rect 189510 150502 189562 150554
rect 189614 150502 189666 150554
rect 189718 150502 204736 150554
rect 1344 150468 204736 150502
rect 1344 149770 204736 149804
rect 1344 149718 4478 149770
rect 4530 149718 4582 149770
rect 4634 149718 4686 149770
rect 4738 149718 35198 149770
rect 35250 149718 35302 149770
rect 35354 149718 35406 149770
rect 35458 149718 65918 149770
rect 65970 149718 66022 149770
rect 66074 149718 66126 149770
rect 66178 149718 96638 149770
rect 96690 149718 96742 149770
rect 96794 149718 96846 149770
rect 96898 149718 127358 149770
rect 127410 149718 127462 149770
rect 127514 149718 127566 149770
rect 127618 149718 158078 149770
rect 158130 149718 158182 149770
rect 158234 149718 158286 149770
rect 158338 149718 188798 149770
rect 188850 149718 188902 149770
rect 188954 149718 189006 149770
rect 189058 149718 204736 149770
rect 1344 149684 204736 149718
rect 1344 148986 204736 149020
rect 1344 148934 5138 148986
rect 5190 148934 5242 148986
rect 5294 148934 5346 148986
rect 5398 148934 35858 148986
rect 35910 148934 35962 148986
rect 36014 148934 36066 148986
rect 36118 148934 66578 148986
rect 66630 148934 66682 148986
rect 66734 148934 66786 148986
rect 66838 148934 97298 148986
rect 97350 148934 97402 148986
rect 97454 148934 97506 148986
rect 97558 148934 128018 148986
rect 128070 148934 128122 148986
rect 128174 148934 128226 148986
rect 128278 148934 158738 148986
rect 158790 148934 158842 148986
rect 158894 148934 158946 148986
rect 158998 148934 189458 148986
rect 189510 148934 189562 148986
rect 189614 148934 189666 148986
rect 189718 148934 204736 148986
rect 1344 148900 204736 148934
rect 1344 148202 204736 148236
rect 1344 148150 4478 148202
rect 4530 148150 4582 148202
rect 4634 148150 4686 148202
rect 4738 148150 35198 148202
rect 35250 148150 35302 148202
rect 35354 148150 35406 148202
rect 35458 148150 65918 148202
rect 65970 148150 66022 148202
rect 66074 148150 66126 148202
rect 66178 148150 96638 148202
rect 96690 148150 96742 148202
rect 96794 148150 96846 148202
rect 96898 148150 127358 148202
rect 127410 148150 127462 148202
rect 127514 148150 127566 148202
rect 127618 148150 158078 148202
rect 158130 148150 158182 148202
rect 158234 148150 158286 148202
rect 158338 148150 188798 148202
rect 188850 148150 188902 148202
rect 188954 148150 189006 148202
rect 189058 148150 204736 148202
rect 1344 148116 204736 148150
rect 1344 147418 204736 147452
rect 1344 147366 5138 147418
rect 5190 147366 5242 147418
rect 5294 147366 5346 147418
rect 5398 147366 35858 147418
rect 35910 147366 35962 147418
rect 36014 147366 36066 147418
rect 36118 147366 66578 147418
rect 66630 147366 66682 147418
rect 66734 147366 66786 147418
rect 66838 147366 97298 147418
rect 97350 147366 97402 147418
rect 97454 147366 97506 147418
rect 97558 147366 128018 147418
rect 128070 147366 128122 147418
rect 128174 147366 128226 147418
rect 128278 147366 158738 147418
rect 158790 147366 158842 147418
rect 158894 147366 158946 147418
rect 158998 147366 189458 147418
rect 189510 147366 189562 147418
rect 189614 147366 189666 147418
rect 189718 147366 204736 147418
rect 1344 147332 204736 147366
rect 1810 146974 1822 147026
rect 1874 146974 1886 147026
rect 2818 146862 2830 146914
rect 2882 146862 2894 146914
rect 1344 146634 204736 146668
rect 1344 146582 4478 146634
rect 4530 146582 4582 146634
rect 4634 146582 4686 146634
rect 4738 146582 35198 146634
rect 35250 146582 35302 146634
rect 35354 146582 35406 146634
rect 35458 146582 65918 146634
rect 65970 146582 66022 146634
rect 66074 146582 66126 146634
rect 66178 146582 96638 146634
rect 96690 146582 96742 146634
rect 96794 146582 96846 146634
rect 96898 146582 127358 146634
rect 127410 146582 127462 146634
rect 127514 146582 127566 146634
rect 127618 146582 158078 146634
rect 158130 146582 158182 146634
rect 158234 146582 158286 146634
rect 158338 146582 188798 146634
rect 188850 146582 188902 146634
rect 188954 146582 189006 146634
rect 189058 146582 204736 146634
rect 1344 146548 204736 146582
rect 1822 146354 1874 146366
rect 1822 146290 1874 146302
rect 204094 146354 204146 146366
rect 204094 146290 204146 146302
rect 201070 146242 201122 146254
rect 201730 146190 201742 146242
rect 201794 146190 201806 146242
rect 201070 146178 201122 146190
rect 1344 145850 204736 145884
rect 1344 145798 5138 145850
rect 5190 145798 5242 145850
rect 5294 145798 5346 145850
rect 5398 145798 35858 145850
rect 35910 145798 35962 145850
rect 36014 145798 36066 145850
rect 36118 145798 66578 145850
rect 66630 145798 66682 145850
rect 66734 145798 66786 145850
rect 66838 145798 97298 145850
rect 97350 145798 97402 145850
rect 97454 145798 97506 145850
rect 97558 145798 128018 145850
rect 128070 145798 128122 145850
rect 128174 145798 128226 145850
rect 128278 145798 158738 145850
rect 158790 145798 158842 145850
rect 158894 145798 158946 145850
rect 158998 145798 189458 145850
rect 189510 145798 189562 145850
rect 189614 145798 189666 145850
rect 189718 145798 204736 145850
rect 1344 145764 204736 145798
rect 1344 145066 204736 145100
rect 1344 145014 4478 145066
rect 4530 145014 4582 145066
rect 4634 145014 4686 145066
rect 4738 145014 35198 145066
rect 35250 145014 35302 145066
rect 35354 145014 35406 145066
rect 35458 145014 65918 145066
rect 65970 145014 66022 145066
rect 66074 145014 66126 145066
rect 66178 145014 96638 145066
rect 96690 145014 96742 145066
rect 96794 145014 96846 145066
rect 96898 145014 127358 145066
rect 127410 145014 127462 145066
rect 127514 145014 127566 145066
rect 127618 145014 158078 145066
rect 158130 145014 158182 145066
rect 158234 145014 158286 145066
rect 158338 145014 188798 145066
rect 188850 145014 188902 145066
rect 188954 145014 189006 145066
rect 189058 145014 204736 145066
rect 1344 144980 204736 145014
rect 1344 144282 17920 144316
rect 1344 144230 5138 144282
rect 5190 144230 5242 144282
rect 5294 144230 5346 144282
rect 5398 144230 17920 144282
rect 1344 144196 17920 144230
rect 188272 144282 204736 144316
rect 188272 144230 189458 144282
rect 189510 144230 189562 144282
rect 189614 144230 189666 144282
rect 189718 144230 204736 144282
rect 188272 144196 204736 144230
rect 1344 143498 17920 143532
rect 1344 143446 4478 143498
rect 4530 143446 4582 143498
rect 4634 143446 4686 143498
rect 4738 143446 17920 143498
rect 1344 143412 17920 143446
rect 188272 143498 204736 143532
rect 188272 143446 188798 143498
rect 188850 143446 188902 143498
rect 188954 143446 189006 143498
rect 189058 143446 204736 143498
rect 188272 143412 204736 143446
rect 1710 142882 1762 142894
rect 1710 142818 1762 142830
rect 1344 142714 17920 142748
rect 1344 142662 5138 142714
rect 5190 142662 5242 142714
rect 5294 142662 5346 142714
rect 5398 142662 17920 142714
rect 1344 142628 17920 142662
rect 188272 142714 204736 142748
rect 188272 142662 189458 142714
rect 189510 142662 189562 142714
rect 189614 142662 189666 142714
rect 189718 142662 204736 142714
rect 188272 142628 204736 142662
rect 1344 141930 17920 141964
rect 1344 141878 4478 141930
rect 4530 141878 4582 141930
rect 4634 141878 4686 141930
rect 4738 141878 17920 141930
rect 1344 141844 17920 141878
rect 188272 141930 204736 141964
rect 188272 141878 188798 141930
rect 188850 141878 188902 141930
rect 188954 141878 189006 141930
rect 189058 141878 204736 141930
rect 188272 141844 204736 141878
rect 1344 141146 17920 141180
rect 1344 141094 5138 141146
rect 5190 141094 5242 141146
rect 5294 141094 5346 141146
rect 5398 141094 17920 141146
rect 1344 141060 17920 141094
rect 188272 141146 204736 141180
rect 188272 141094 189458 141146
rect 189510 141094 189562 141146
rect 189614 141094 189666 141146
rect 189718 141094 204736 141146
rect 188272 141060 204736 141094
rect 1344 140362 17920 140396
rect 1344 140310 4478 140362
rect 4530 140310 4582 140362
rect 4634 140310 4686 140362
rect 4738 140310 17920 140362
rect 1344 140276 17920 140310
rect 188272 140362 204736 140396
rect 188272 140310 188798 140362
rect 188850 140310 188902 140362
rect 188954 140310 189006 140362
rect 189058 140310 204736 140362
rect 188272 140276 204736 140310
rect 1344 139578 17920 139612
rect 1344 139526 5138 139578
rect 5190 139526 5242 139578
rect 5294 139526 5346 139578
rect 5398 139526 17920 139578
rect 1344 139492 17920 139526
rect 188272 139578 204736 139612
rect 188272 139526 189458 139578
rect 189510 139526 189562 139578
rect 189614 139526 189666 139578
rect 189718 139526 204736 139578
rect 188272 139492 204736 139526
rect 1710 138962 1762 138974
rect 1710 138898 1762 138910
rect 1344 138794 17920 138828
rect 1344 138742 4478 138794
rect 4530 138742 4582 138794
rect 4634 138742 4686 138794
rect 4738 138742 17920 138794
rect 1344 138708 17920 138742
rect 188272 138794 204736 138828
rect 188272 138742 188798 138794
rect 188850 138742 188902 138794
rect 188954 138742 189006 138794
rect 189058 138742 204736 138794
rect 188272 138708 204736 138742
rect 1344 138010 17920 138044
rect 1344 137958 5138 138010
rect 5190 137958 5242 138010
rect 5294 137958 5346 138010
rect 5398 137958 17920 138010
rect 1344 137924 17920 137958
rect 188272 138010 204736 138044
rect 188272 137958 189458 138010
rect 189510 137958 189562 138010
rect 189614 137958 189666 138010
rect 189718 137958 204736 138010
rect 188272 137924 204736 137958
rect 1344 137226 17920 137260
rect 1344 137174 4478 137226
rect 4530 137174 4582 137226
rect 4634 137174 4686 137226
rect 4738 137174 17920 137226
rect 1344 137140 17920 137174
rect 188272 137226 204736 137260
rect 188272 137174 188798 137226
rect 188850 137174 188902 137226
rect 188954 137174 189006 137226
rect 189058 137174 204736 137226
rect 188272 137140 204736 137174
rect 1344 136442 17920 136476
rect 1344 136390 5138 136442
rect 5190 136390 5242 136442
rect 5294 136390 5346 136442
rect 5398 136390 17920 136442
rect 1344 136356 17920 136390
rect 188272 136442 204736 136476
rect 188272 136390 189458 136442
rect 189510 136390 189562 136442
rect 189614 136390 189666 136442
rect 189718 136390 204736 136442
rect 188272 136356 204736 136390
rect 1344 135658 17920 135692
rect 1344 135606 4478 135658
rect 4530 135606 4582 135658
rect 4634 135606 4686 135658
rect 4738 135606 17920 135658
rect 1344 135572 17920 135606
rect 188272 135658 204736 135692
rect 188272 135606 188798 135658
rect 188850 135606 188902 135658
rect 188954 135606 189006 135658
rect 189058 135606 204736 135658
rect 188272 135572 204736 135606
rect 1698 135214 1710 135266
rect 1762 135214 1774 135266
rect 2818 135102 2830 135154
rect 2882 135102 2894 135154
rect 1344 134874 17920 134908
rect 1344 134822 5138 134874
rect 5190 134822 5242 134874
rect 5294 134822 5346 134874
rect 5398 134822 17920 134874
rect 1344 134788 17920 134822
rect 188272 134874 204736 134908
rect 188272 134822 189458 134874
rect 189510 134822 189562 134874
rect 189614 134822 189666 134874
rect 189718 134822 204736 134874
rect 188272 134788 204736 134822
rect 1822 134706 1874 134718
rect 1822 134642 1874 134654
rect 1344 134090 17920 134124
rect 1344 134038 4478 134090
rect 4530 134038 4582 134090
rect 4634 134038 4686 134090
rect 4738 134038 17920 134090
rect 1344 134004 17920 134038
rect 188272 134090 204736 134124
rect 188272 134038 188798 134090
rect 188850 134038 188902 134090
rect 188954 134038 189006 134090
rect 189058 134038 204736 134090
rect 188272 134004 204736 134038
rect 1344 133306 17920 133340
rect 1344 133254 5138 133306
rect 5190 133254 5242 133306
rect 5294 133254 5346 133306
rect 5398 133254 17920 133306
rect 1344 133220 17920 133254
rect 188272 133306 204736 133340
rect 188272 133254 189458 133306
rect 189510 133254 189562 133306
rect 189614 133254 189666 133306
rect 189718 133254 204736 133306
rect 188272 133220 204736 133254
rect 1344 132522 17920 132556
rect 1344 132470 4478 132522
rect 4530 132470 4582 132522
rect 4634 132470 4686 132522
rect 4738 132470 17920 132522
rect 1344 132436 17920 132470
rect 188272 132522 204736 132556
rect 188272 132470 188798 132522
rect 188850 132470 188902 132522
rect 188954 132470 189006 132522
rect 189058 132470 204736 132522
rect 188272 132436 204736 132470
rect 1710 131906 1762 131918
rect 1710 131842 1762 131854
rect 1344 131738 17920 131772
rect 1344 131686 5138 131738
rect 5190 131686 5242 131738
rect 5294 131686 5346 131738
rect 5398 131686 17920 131738
rect 1344 131652 17920 131686
rect 188272 131738 204736 131772
rect 188272 131686 189458 131738
rect 189510 131686 189562 131738
rect 189614 131686 189666 131738
rect 189718 131686 204736 131738
rect 188272 131652 204736 131686
rect 1344 130954 17920 130988
rect 1344 130902 4478 130954
rect 4530 130902 4582 130954
rect 4634 130902 4686 130954
rect 4738 130902 17920 130954
rect 1344 130868 17920 130902
rect 188272 130954 204736 130988
rect 188272 130902 188798 130954
rect 188850 130902 188902 130954
rect 188954 130902 189006 130954
rect 189058 130902 204736 130954
rect 188272 130868 204736 130902
rect 1344 130170 17920 130204
rect 1344 130118 5138 130170
rect 5190 130118 5242 130170
rect 5294 130118 5346 130170
rect 5398 130118 17920 130170
rect 1344 130084 17920 130118
rect 188272 130170 204736 130204
rect 188272 130118 189458 130170
rect 189510 130118 189562 130170
rect 189614 130118 189666 130170
rect 189718 130118 204736 130170
rect 188272 130084 204736 130118
rect 1344 129386 17920 129420
rect 1344 129334 4478 129386
rect 4530 129334 4582 129386
rect 4634 129334 4686 129386
rect 4738 129334 17920 129386
rect 1344 129300 17920 129334
rect 188272 129386 204736 129420
rect 188272 129334 188798 129386
rect 188850 129334 188902 129386
rect 188954 129334 189006 129386
rect 189058 129334 204736 129386
rect 188272 129300 204736 129334
rect 1344 128602 17920 128636
rect 1344 128550 5138 128602
rect 5190 128550 5242 128602
rect 5294 128550 5346 128602
rect 5398 128550 17920 128602
rect 1344 128516 17920 128550
rect 188272 128602 204736 128636
rect 188272 128550 189458 128602
rect 189510 128550 189562 128602
rect 189614 128550 189666 128602
rect 189718 128550 204736 128602
rect 188272 128516 204736 128550
rect 203758 128322 203810 128334
rect 203758 128258 203810 128270
rect 1710 127986 1762 127998
rect 1710 127922 1762 127934
rect 1344 127818 17920 127852
rect 1344 127766 4478 127818
rect 4530 127766 4582 127818
rect 4634 127766 4686 127818
rect 4738 127766 17920 127818
rect 1344 127732 17920 127766
rect 188272 127818 204736 127852
rect 188272 127766 188798 127818
rect 188850 127766 188902 127818
rect 188954 127766 189006 127818
rect 189058 127766 204736 127818
rect 188272 127732 204736 127766
rect 1344 127034 17920 127068
rect 1344 126982 5138 127034
rect 5190 126982 5242 127034
rect 5294 126982 5346 127034
rect 5398 126982 17920 127034
rect 1344 126948 17920 126982
rect 188272 127034 204736 127068
rect 188272 126982 189458 127034
rect 189510 126982 189562 127034
rect 189614 126982 189666 127034
rect 189718 126982 204736 127034
rect 188272 126948 204736 126982
rect 1344 126250 17920 126284
rect 1344 126198 4478 126250
rect 4530 126198 4582 126250
rect 4634 126198 4686 126250
rect 4738 126198 17920 126250
rect 1344 126164 17920 126198
rect 188272 126250 204736 126284
rect 188272 126198 188798 126250
rect 188850 126198 188902 126250
rect 188954 126198 189006 126250
rect 189058 126198 204736 126250
rect 188272 126164 204736 126198
rect 1344 125466 17920 125500
rect 1344 125414 5138 125466
rect 5190 125414 5242 125466
rect 5294 125414 5346 125466
rect 5398 125414 17920 125466
rect 1344 125380 17920 125414
rect 188272 125466 204736 125500
rect 188272 125414 189458 125466
rect 189510 125414 189562 125466
rect 189614 125414 189666 125466
rect 189718 125414 204736 125466
rect 188272 125380 204736 125414
rect 1344 124682 17920 124716
rect 1344 124630 4478 124682
rect 4530 124630 4582 124682
rect 4634 124630 4686 124682
rect 4738 124630 17920 124682
rect 1344 124596 17920 124630
rect 188272 124682 204736 124716
rect 188272 124630 188798 124682
rect 188850 124630 188902 124682
rect 188954 124630 189006 124682
rect 189058 124630 204736 124682
rect 188272 124596 204736 124630
rect 1810 124238 1822 124290
rect 1874 124238 1886 124290
rect 2818 124126 2830 124178
rect 2882 124126 2894 124178
rect 1344 123898 17920 123932
rect 1344 123846 5138 123898
rect 5190 123846 5242 123898
rect 5294 123846 5346 123898
rect 5398 123846 17920 123898
rect 1344 123812 17920 123846
rect 188272 123898 204736 123932
rect 188272 123846 189458 123898
rect 189510 123846 189562 123898
rect 189614 123846 189666 123898
rect 189718 123846 204736 123898
rect 188272 123812 204736 123846
rect 1822 123730 1874 123742
rect 1822 123666 1874 123678
rect 1344 123114 17920 123148
rect 1344 123062 4478 123114
rect 4530 123062 4582 123114
rect 4634 123062 4686 123114
rect 4738 123062 17920 123114
rect 1344 123028 17920 123062
rect 188272 123114 204736 123148
rect 188272 123062 188798 123114
rect 188850 123062 188902 123114
rect 188954 123062 189006 123114
rect 189058 123062 204736 123114
rect 188272 123028 204736 123062
rect 1344 122330 17920 122364
rect 1344 122278 5138 122330
rect 5190 122278 5242 122330
rect 5294 122278 5346 122330
rect 5398 122278 17920 122330
rect 1344 122244 17920 122278
rect 188272 122330 204736 122364
rect 188272 122278 189458 122330
rect 189510 122278 189562 122330
rect 189614 122278 189666 122330
rect 189718 122278 204736 122330
rect 188272 122244 204736 122278
rect 1344 121546 17920 121580
rect 1344 121494 4478 121546
rect 4530 121494 4582 121546
rect 4634 121494 4686 121546
rect 4738 121494 17920 121546
rect 1344 121460 17920 121494
rect 188272 121546 204736 121580
rect 188272 121494 188798 121546
rect 188850 121494 188902 121546
rect 188954 121494 189006 121546
rect 189058 121494 204736 121546
rect 188272 121460 204736 121494
rect 1344 120762 17920 120796
rect 1344 120710 5138 120762
rect 5190 120710 5242 120762
rect 5294 120710 5346 120762
rect 5398 120710 17920 120762
rect 1344 120676 17920 120710
rect 188272 120762 204736 120796
rect 188272 120710 189458 120762
rect 189510 120710 189562 120762
rect 189614 120710 189666 120762
rect 189718 120710 204736 120762
rect 188272 120676 204736 120710
rect 1710 120482 1762 120494
rect 1710 120418 1762 120430
rect 1344 119978 17920 120012
rect 1344 119926 4478 119978
rect 4530 119926 4582 119978
rect 4634 119926 4686 119978
rect 4738 119926 17920 119978
rect 1344 119892 17920 119926
rect 188272 119978 204736 120012
rect 188272 119926 188798 119978
rect 188850 119926 188902 119978
rect 188954 119926 189006 119978
rect 189058 119926 204736 119978
rect 188272 119892 204736 119926
rect 204094 119698 204146 119710
rect 204094 119634 204146 119646
rect 202178 119534 202190 119586
rect 202242 119534 202254 119586
rect 1344 119194 17920 119228
rect 1344 119142 5138 119194
rect 5190 119142 5242 119194
rect 5294 119142 5346 119194
rect 5398 119142 17920 119194
rect 1344 119108 17920 119142
rect 188272 119194 204736 119228
rect 188272 119142 189458 119194
rect 189510 119142 189562 119194
rect 189614 119142 189666 119194
rect 189718 119142 204736 119194
rect 188272 119108 204736 119142
rect 203758 118690 203810 118702
rect 203758 118626 203810 118638
rect 1344 118410 17920 118444
rect 1344 118358 4478 118410
rect 4530 118358 4582 118410
rect 4634 118358 4686 118410
rect 4738 118358 17920 118410
rect 1344 118324 17920 118358
rect 188272 118410 204736 118444
rect 188272 118358 188798 118410
rect 188850 118358 188902 118410
rect 188954 118358 189006 118410
rect 189058 118358 204736 118410
rect 188272 118324 204736 118358
rect 1344 117626 17920 117660
rect 1344 117574 5138 117626
rect 5190 117574 5242 117626
rect 5294 117574 5346 117626
rect 5398 117574 17920 117626
rect 1344 117540 17920 117574
rect 188272 117626 204736 117660
rect 188272 117574 189458 117626
rect 189510 117574 189562 117626
rect 189614 117574 189666 117626
rect 189718 117574 204736 117626
rect 188272 117540 204736 117574
rect 1344 116842 17920 116876
rect 1344 116790 4478 116842
rect 4530 116790 4582 116842
rect 4634 116790 4686 116842
rect 4738 116790 17920 116842
rect 1344 116756 17920 116790
rect 188272 116842 204736 116876
rect 188272 116790 188798 116842
rect 188850 116790 188902 116842
rect 188954 116790 189006 116842
rect 189058 116790 204736 116842
rect 188272 116756 204736 116790
rect 1710 116562 1762 116574
rect 1710 116498 1762 116510
rect 1344 116058 17920 116092
rect 1344 116006 5138 116058
rect 5190 116006 5242 116058
rect 5294 116006 5346 116058
rect 5398 116006 17920 116058
rect 1344 115972 17920 116006
rect 188272 116058 204736 116092
rect 188272 116006 189458 116058
rect 189510 116006 189562 116058
rect 189614 116006 189666 116058
rect 189718 116006 204736 116058
rect 188272 115972 204736 116006
rect 1344 115274 17920 115308
rect 1344 115222 4478 115274
rect 4530 115222 4582 115274
rect 4634 115222 4686 115274
rect 4738 115222 17920 115274
rect 1344 115188 17920 115222
rect 188272 115274 204736 115308
rect 188272 115222 188798 115274
rect 188850 115222 188902 115274
rect 188954 115222 189006 115274
rect 189058 115222 204736 115274
rect 188272 115188 204736 115222
rect 1344 114490 17920 114524
rect 1344 114438 5138 114490
rect 5190 114438 5242 114490
rect 5294 114438 5346 114490
rect 5398 114438 17920 114490
rect 1344 114404 17920 114438
rect 188272 114490 204736 114524
rect 188272 114438 189458 114490
rect 189510 114438 189562 114490
rect 189614 114438 189666 114490
rect 189718 114438 204736 114490
rect 188272 114404 204736 114438
rect 1344 113706 17920 113740
rect 1344 113654 4478 113706
rect 4530 113654 4582 113706
rect 4634 113654 4686 113706
rect 4738 113654 17920 113706
rect 1344 113620 17920 113654
rect 188272 113706 204736 113740
rect 188272 113654 188798 113706
rect 188850 113654 188902 113706
rect 188954 113654 189006 113706
rect 189058 113654 204736 113706
rect 188272 113620 204736 113654
rect 1344 112922 17920 112956
rect 1344 112870 5138 112922
rect 5190 112870 5242 112922
rect 5294 112870 5346 112922
rect 5398 112870 17920 112922
rect 1344 112836 17920 112870
rect 188272 112922 204736 112956
rect 188272 112870 189458 112922
rect 189510 112870 189562 112922
rect 189614 112870 189666 112922
rect 189718 112870 204736 112922
rect 188272 112836 204736 112870
rect 1698 112478 1710 112530
rect 1762 112478 1774 112530
rect 2818 112366 2830 112418
rect 2882 112366 2894 112418
rect 1344 112138 17920 112172
rect 1344 112086 4478 112138
rect 4530 112086 4582 112138
rect 4634 112086 4686 112138
rect 4738 112086 17920 112138
rect 1344 112052 17920 112086
rect 188272 112138 204736 112172
rect 188272 112086 188798 112138
rect 188850 112086 188902 112138
rect 188954 112086 189006 112138
rect 189058 112086 204736 112138
rect 188272 112052 204736 112086
rect 1822 111858 1874 111870
rect 1822 111794 1874 111806
rect 1344 111354 17920 111388
rect 1344 111302 5138 111354
rect 5190 111302 5242 111354
rect 5294 111302 5346 111354
rect 5398 111302 17920 111354
rect 1344 111268 17920 111302
rect 188272 111354 204736 111388
rect 188272 111302 189458 111354
rect 189510 111302 189562 111354
rect 189614 111302 189666 111354
rect 189718 111302 204736 111354
rect 188272 111268 204736 111302
rect 1344 110570 17920 110604
rect 1344 110518 4478 110570
rect 4530 110518 4582 110570
rect 4634 110518 4686 110570
rect 4738 110518 17920 110570
rect 1344 110484 17920 110518
rect 188272 110570 204736 110604
rect 188272 110518 188798 110570
rect 188850 110518 188902 110570
rect 188954 110518 189006 110570
rect 189058 110518 204736 110570
rect 188272 110484 204736 110518
rect 1344 109786 17920 109820
rect 1344 109734 5138 109786
rect 5190 109734 5242 109786
rect 5294 109734 5346 109786
rect 5398 109734 17920 109786
rect 1344 109700 17920 109734
rect 188272 109786 204736 109820
rect 188272 109734 189458 109786
rect 189510 109734 189562 109786
rect 189614 109734 189666 109786
rect 189718 109734 204736 109786
rect 188272 109700 204736 109734
rect 1344 109002 17920 109036
rect 1344 108950 4478 109002
rect 4530 108950 4582 109002
rect 4634 108950 4686 109002
rect 4738 108950 17920 109002
rect 1344 108916 17920 108950
rect 188272 109002 204736 109036
rect 188272 108950 188798 109002
rect 188850 108950 188902 109002
rect 188954 108950 189006 109002
rect 189058 108950 204736 109002
rect 188272 108916 204736 108950
rect 1710 108498 1762 108510
rect 1710 108434 1762 108446
rect 1344 108218 17920 108252
rect 1344 108166 5138 108218
rect 5190 108166 5242 108218
rect 5294 108166 5346 108218
rect 5398 108166 17920 108218
rect 1344 108132 17920 108166
rect 188272 108218 204736 108252
rect 188272 108166 189458 108218
rect 189510 108166 189562 108218
rect 189614 108166 189666 108218
rect 189718 108166 204736 108218
rect 188272 108132 204736 108166
rect 1344 107434 17920 107468
rect 1344 107382 4478 107434
rect 4530 107382 4582 107434
rect 4634 107382 4686 107434
rect 4738 107382 17920 107434
rect 1344 107348 17920 107382
rect 188272 107434 204736 107468
rect 188272 107382 188798 107434
rect 188850 107382 188902 107434
rect 188954 107382 189006 107434
rect 189058 107382 204736 107434
rect 188272 107348 204736 107382
rect 1344 106650 17920 106684
rect 1344 106598 5138 106650
rect 5190 106598 5242 106650
rect 5294 106598 5346 106650
rect 5398 106598 17920 106650
rect 1344 106564 17920 106598
rect 188272 106650 204736 106684
rect 188272 106598 189458 106650
rect 189510 106598 189562 106650
rect 189614 106598 189666 106650
rect 189718 106598 204736 106650
rect 188272 106564 204736 106598
rect 1344 105866 17920 105900
rect 1344 105814 4478 105866
rect 4530 105814 4582 105866
rect 4634 105814 4686 105866
rect 4738 105814 17920 105866
rect 1344 105780 17920 105814
rect 188272 105866 204736 105900
rect 188272 105814 188798 105866
rect 188850 105814 188902 105866
rect 188954 105814 189006 105866
rect 189058 105814 204736 105866
rect 188272 105780 204736 105814
rect 1710 105586 1762 105598
rect 1710 105522 1762 105534
rect 1344 105082 17920 105116
rect 1344 105030 5138 105082
rect 5190 105030 5242 105082
rect 5294 105030 5346 105082
rect 5398 105030 17920 105082
rect 1344 104996 17920 105030
rect 188272 105082 204736 105116
rect 188272 105030 189458 105082
rect 189510 105030 189562 105082
rect 189614 105030 189666 105082
rect 189718 105030 204736 105082
rect 188272 104996 204736 105030
rect 1344 104298 17920 104332
rect 1344 104246 4478 104298
rect 4530 104246 4582 104298
rect 4634 104246 4686 104298
rect 4738 104246 17920 104298
rect 1344 104212 17920 104246
rect 188272 104298 204736 104332
rect 188272 104246 188798 104298
rect 188850 104246 188902 104298
rect 188954 104246 189006 104298
rect 189058 104246 204736 104298
rect 188272 104212 204736 104246
rect 1344 103514 17920 103548
rect 1344 103462 5138 103514
rect 5190 103462 5242 103514
rect 5294 103462 5346 103514
rect 5398 103462 17920 103514
rect 1344 103428 17920 103462
rect 188272 103514 204736 103548
rect 188272 103462 189458 103514
rect 189510 103462 189562 103514
rect 189614 103462 189666 103514
rect 189718 103462 204736 103514
rect 188272 103428 204736 103462
rect 1344 102730 17920 102764
rect 1344 102678 4478 102730
rect 4530 102678 4582 102730
rect 4634 102678 4686 102730
rect 4738 102678 17920 102730
rect 1344 102644 17920 102678
rect 188272 102730 204736 102764
rect 188272 102678 188798 102730
rect 188850 102678 188902 102730
rect 188954 102678 189006 102730
rect 189058 102678 204736 102730
rect 188272 102644 204736 102678
rect 204318 102114 204370 102126
rect 204318 102050 204370 102062
rect 1344 101946 17920 101980
rect 1344 101894 5138 101946
rect 5190 101894 5242 101946
rect 5294 101894 5346 101946
rect 5398 101894 17920 101946
rect 1344 101860 17920 101894
rect 188272 101946 204736 101980
rect 188272 101894 189458 101946
rect 189510 101894 189562 101946
rect 189614 101894 189666 101946
rect 189718 101894 204736 101946
rect 188272 101860 204736 101894
rect 2034 101614 2046 101666
rect 2098 101614 2110 101666
rect 1710 101554 1762 101566
rect 1710 101490 1762 101502
rect 2494 101442 2546 101454
rect 2494 101378 2546 101390
rect 1344 101162 17920 101196
rect 1344 101110 4478 101162
rect 4530 101110 4582 101162
rect 4634 101110 4686 101162
rect 4738 101110 17920 101162
rect 1344 101076 17920 101110
rect 188272 101162 204736 101196
rect 188272 101110 188798 101162
rect 188850 101110 188902 101162
rect 188954 101110 189006 101162
rect 189058 101110 204736 101162
rect 188272 101076 204736 101110
rect 1344 100378 17920 100412
rect 1344 100326 5138 100378
rect 5190 100326 5242 100378
rect 5294 100326 5346 100378
rect 5398 100326 17920 100378
rect 1344 100292 17920 100326
rect 188272 100378 204736 100412
rect 188272 100326 189458 100378
rect 189510 100326 189562 100378
rect 189614 100326 189666 100378
rect 189718 100326 204736 100378
rect 188272 100292 204736 100326
rect 1344 99594 17920 99628
rect 1344 99542 4478 99594
rect 4530 99542 4582 99594
rect 4634 99542 4686 99594
rect 4738 99542 17920 99594
rect 1344 99508 17920 99542
rect 188272 99594 204736 99628
rect 188272 99542 188798 99594
rect 188850 99542 188902 99594
rect 188954 99542 189006 99594
rect 189058 99542 204736 99594
rect 188272 99508 204736 99542
rect 1344 98810 17920 98844
rect 1344 98758 5138 98810
rect 5190 98758 5242 98810
rect 5294 98758 5346 98810
rect 5398 98758 17920 98810
rect 1344 98724 17920 98758
rect 188272 98810 204736 98844
rect 188272 98758 189458 98810
rect 189510 98758 189562 98810
rect 189614 98758 189666 98810
rect 189718 98758 204736 98810
rect 188272 98724 204736 98758
rect 1344 98026 17920 98060
rect 1344 97974 4478 98026
rect 4530 97974 4582 98026
rect 4634 97974 4686 98026
rect 4738 97974 17920 98026
rect 1344 97940 17920 97974
rect 188272 98026 204736 98060
rect 188272 97974 188798 98026
rect 188850 97974 188902 98026
rect 188954 97974 189006 98026
rect 189058 97974 204736 98026
rect 188272 97940 204736 97974
rect 1710 97410 1762 97422
rect 1710 97346 1762 97358
rect 1344 97242 17920 97276
rect 1344 97190 5138 97242
rect 5190 97190 5242 97242
rect 5294 97190 5346 97242
rect 5398 97190 17920 97242
rect 1344 97156 17920 97190
rect 188272 97242 204736 97276
rect 188272 97190 189458 97242
rect 189510 97190 189562 97242
rect 189614 97190 189666 97242
rect 189718 97190 204736 97242
rect 188272 97156 204736 97190
rect 1344 96458 17920 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 17920 96458
rect 1344 96372 17920 96406
rect 188272 96458 204736 96492
rect 188272 96406 188798 96458
rect 188850 96406 188902 96458
rect 188954 96406 189006 96458
rect 189058 96406 204736 96458
rect 188272 96372 204736 96406
rect 1344 95674 17920 95708
rect 1344 95622 5138 95674
rect 5190 95622 5242 95674
rect 5294 95622 5346 95674
rect 5398 95622 17920 95674
rect 1344 95588 17920 95622
rect 188272 95674 204736 95708
rect 188272 95622 189458 95674
rect 189510 95622 189562 95674
rect 189614 95622 189666 95674
rect 189718 95622 204736 95674
rect 188272 95588 204736 95622
rect 1344 94890 17920 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 17920 94890
rect 1344 94804 17920 94838
rect 188272 94890 204736 94924
rect 188272 94838 188798 94890
rect 188850 94838 188902 94890
rect 188954 94838 189006 94890
rect 189058 94838 204736 94890
rect 188272 94804 204736 94838
rect 1344 94106 17920 94140
rect 1344 94054 5138 94106
rect 5190 94054 5242 94106
rect 5294 94054 5346 94106
rect 5398 94054 17920 94106
rect 1344 94020 17920 94054
rect 188272 94106 204736 94140
rect 188272 94054 189458 94106
rect 189510 94054 189562 94106
rect 189614 94054 189666 94106
rect 189718 94054 204736 94106
rect 188272 94020 204736 94054
rect 201170 93662 201182 93714
rect 201234 93662 201246 93714
rect 203186 93550 203198 93602
rect 203250 93550 203262 93602
rect 1710 93490 1762 93502
rect 1710 93426 1762 93438
rect 1344 93322 17920 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 17920 93322
rect 1344 93236 17920 93270
rect 188272 93322 204736 93356
rect 188272 93270 188798 93322
rect 188850 93270 188902 93322
rect 188954 93270 189006 93322
rect 189058 93270 204736 93322
rect 188272 93236 204736 93270
rect 203982 93042 204034 93054
rect 203982 92978 204034 92990
rect 1344 92538 17920 92572
rect 1344 92486 5138 92538
rect 5190 92486 5242 92538
rect 5294 92486 5346 92538
rect 5398 92486 17920 92538
rect 1344 92452 17920 92486
rect 188272 92538 204736 92572
rect 188272 92486 189458 92538
rect 189510 92486 189562 92538
rect 189614 92486 189666 92538
rect 189718 92486 204736 92538
rect 188272 92452 204736 92486
rect 1344 91754 17920 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 17920 91754
rect 1344 91668 17920 91702
rect 188272 91754 204736 91788
rect 188272 91702 188798 91754
rect 188850 91702 188902 91754
rect 188954 91702 189006 91754
rect 189058 91702 204736 91754
rect 188272 91668 204736 91702
rect 1344 90970 17920 91004
rect 1344 90918 5138 90970
rect 5190 90918 5242 90970
rect 5294 90918 5346 90970
rect 5398 90918 17920 90970
rect 1344 90884 17920 90918
rect 188272 90970 204736 91004
rect 188272 90918 189458 90970
rect 189510 90918 189562 90970
rect 189614 90918 189666 90970
rect 189718 90918 204736 90970
rect 188272 90884 204736 90918
rect 1344 90186 17920 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 17920 90186
rect 1344 90100 17920 90134
rect 188272 90186 204736 90220
rect 188272 90134 188798 90186
rect 188850 90134 188902 90186
rect 188954 90134 189006 90186
rect 189058 90134 204736 90186
rect 188272 90100 204736 90134
rect 1710 89570 1762 89582
rect 2494 89570 2546 89582
rect 2034 89518 2046 89570
rect 2098 89518 2110 89570
rect 1710 89506 1762 89518
rect 2494 89506 2546 89518
rect 1344 89402 17920 89436
rect 1344 89350 5138 89402
rect 5190 89350 5242 89402
rect 5294 89350 5346 89402
rect 5398 89350 17920 89402
rect 1344 89316 17920 89350
rect 188272 89402 204736 89436
rect 188272 89350 189458 89402
rect 189510 89350 189562 89402
rect 189614 89350 189666 89402
rect 189718 89350 204736 89402
rect 188272 89316 204736 89350
rect 1344 88618 17920 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 17920 88618
rect 1344 88532 17920 88566
rect 188272 88618 204736 88652
rect 188272 88566 188798 88618
rect 188850 88566 188902 88618
rect 188954 88566 189006 88618
rect 189058 88566 204736 88618
rect 188272 88532 204736 88566
rect 1344 87834 17920 87868
rect 1344 87782 5138 87834
rect 5190 87782 5242 87834
rect 5294 87782 5346 87834
rect 5398 87782 17920 87834
rect 1344 87748 17920 87782
rect 188272 87834 204736 87868
rect 188272 87782 189458 87834
rect 189510 87782 189562 87834
rect 189614 87782 189666 87834
rect 189718 87782 204736 87834
rect 188272 87748 204736 87782
rect 1344 87050 17920 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 17920 87050
rect 1344 86964 17920 86998
rect 188272 87050 204736 87084
rect 188272 86998 188798 87050
rect 188850 86998 188902 87050
rect 188954 86998 189006 87050
rect 189058 86998 204736 87050
rect 188272 86964 204736 86998
rect 1344 86266 17920 86300
rect 1344 86214 5138 86266
rect 5190 86214 5242 86266
rect 5294 86214 5346 86266
rect 5398 86214 17920 86266
rect 1344 86180 17920 86214
rect 188272 86266 204736 86300
rect 188272 86214 189458 86266
rect 189510 86214 189562 86266
rect 189614 86214 189666 86266
rect 189718 86214 204736 86266
rect 188272 86180 204736 86214
rect 1710 85986 1762 85998
rect 1710 85922 1762 85934
rect 1344 85482 17920 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 17920 85482
rect 1344 85396 17920 85430
rect 188272 85482 204736 85516
rect 188272 85430 188798 85482
rect 188850 85430 188902 85482
rect 188954 85430 189006 85482
rect 189058 85430 204736 85482
rect 188272 85396 204736 85430
rect 1344 84698 17920 84732
rect 1344 84646 5138 84698
rect 5190 84646 5242 84698
rect 5294 84646 5346 84698
rect 5398 84646 17920 84698
rect 1344 84612 17920 84646
rect 188272 84698 204736 84732
rect 188272 84646 189458 84698
rect 189510 84646 189562 84698
rect 189614 84646 189666 84698
rect 189718 84646 204736 84698
rect 188272 84612 204736 84646
rect 1344 83914 17920 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 17920 83914
rect 1344 83828 17920 83862
rect 188272 83914 204736 83948
rect 188272 83862 188798 83914
rect 188850 83862 188902 83914
rect 188954 83862 189006 83914
rect 189058 83862 204736 83914
rect 188272 83828 204736 83862
rect 1344 83130 17920 83164
rect 1344 83078 5138 83130
rect 5190 83078 5242 83130
rect 5294 83078 5346 83130
rect 5398 83078 17920 83130
rect 1344 83044 17920 83078
rect 188272 83130 204736 83164
rect 188272 83078 189458 83130
rect 189510 83078 189562 83130
rect 189614 83078 189666 83130
rect 189718 83078 204736 83130
rect 188272 83044 204736 83078
rect 1344 82346 17920 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 17920 82346
rect 1344 82260 17920 82294
rect 188272 82346 204736 82380
rect 188272 82294 188798 82346
rect 188850 82294 188902 82346
rect 188954 82294 189006 82346
rect 189058 82294 204736 82346
rect 188272 82260 204736 82294
rect 1710 82066 1762 82078
rect 1710 82002 1762 82014
rect 1344 81562 17920 81596
rect 1344 81510 5138 81562
rect 5190 81510 5242 81562
rect 5294 81510 5346 81562
rect 5398 81510 17920 81562
rect 1344 81476 17920 81510
rect 188272 81562 204736 81596
rect 188272 81510 189458 81562
rect 189510 81510 189562 81562
rect 189614 81510 189666 81562
rect 189718 81510 204736 81562
rect 188272 81476 204736 81510
rect 1344 80778 17920 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 17920 80778
rect 1344 80692 17920 80726
rect 188272 80778 204736 80812
rect 188272 80726 188798 80778
rect 188850 80726 188902 80778
rect 188954 80726 189006 80778
rect 189058 80726 204736 80778
rect 188272 80692 204736 80726
rect 1344 79994 17920 80028
rect 1344 79942 5138 79994
rect 5190 79942 5242 79994
rect 5294 79942 5346 79994
rect 5398 79942 17920 79994
rect 1344 79908 17920 79942
rect 188272 79994 204736 80028
rect 188272 79942 189458 79994
rect 189510 79942 189562 79994
rect 189614 79942 189666 79994
rect 189718 79942 204736 79994
rect 188272 79908 204736 79942
rect 1344 79210 17920 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 17920 79210
rect 1344 79124 17920 79158
rect 188272 79210 204736 79244
rect 188272 79158 188798 79210
rect 188850 79158 188902 79210
rect 188954 79158 189006 79210
rect 189058 79158 204736 79210
rect 188272 79124 204736 79158
rect 1710 78594 1762 78606
rect 2494 78594 2546 78606
rect 2034 78542 2046 78594
rect 2098 78542 2110 78594
rect 1710 78530 1762 78542
rect 2494 78530 2546 78542
rect 17614 78594 17666 78606
rect 17614 78530 17666 78542
rect 1344 78426 17920 78460
rect 1344 78374 5138 78426
rect 5190 78374 5242 78426
rect 5294 78374 5346 78426
rect 5398 78374 17920 78426
rect 1344 78340 17920 78374
rect 188272 78426 204736 78460
rect 188272 78374 189458 78426
rect 189510 78374 189562 78426
rect 189614 78374 189666 78426
rect 189718 78374 204736 78426
rect 188272 78340 204736 78374
rect 17614 77922 17666 77934
rect 17614 77858 17666 77870
rect 1344 77642 17920 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 17920 77642
rect 1344 77556 17920 77590
rect 188272 77642 204736 77676
rect 188272 77590 188798 77642
rect 188850 77590 188902 77642
rect 188954 77590 189006 77642
rect 189058 77590 204736 77642
rect 188272 77556 204736 77590
rect 1344 76858 17920 76892
rect 1344 76806 5138 76858
rect 5190 76806 5242 76858
rect 5294 76806 5346 76858
rect 5398 76806 17920 76858
rect 1344 76772 17920 76806
rect 188272 76858 204736 76892
rect 188272 76806 189458 76858
rect 189510 76806 189562 76858
rect 189614 76806 189666 76858
rect 189718 76806 204736 76858
rect 188272 76772 204736 76806
rect 17614 76354 17666 76366
rect 17614 76290 17666 76302
rect 1344 76074 17920 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 17920 76074
rect 1344 75988 17920 76022
rect 188272 76074 204736 76108
rect 188272 76022 188798 76074
rect 188850 76022 188902 76074
rect 188954 76022 189006 76074
rect 189058 76022 204736 76074
rect 188272 75988 204736 76022
rect 17502 75682 17554 75694
rect 17502 75618 17554 75630
rect 204318 75570 204370 75582
rect 204318 75506 204370 75518
rect 1344 75290 17920 75324
rect 1344 75238 5138 75290
rect 5190 75238 5242 75290
rect 5294 75238 5346 75290
rect 5398 75238 17920 75290
rect 1344 75204 17920 75238
rect 188272 75290 204736 75324
rect 188272 75238 189458 75290
rect 189510 75238 189562 75290
rect 189614 75238 189666 75290
rect 189718 75238 204736 75290
rect 188272 75204 204736 75238
rect 1710 75010 1762 75022
rect 1710 74946 1762 74958
rect 17502 74786 17554 74798
rect 17502 74722 17554 74734
rect 1344 74506 17920 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 17920 74506
rect 1344 74420 17920 74454
rect 188272 74506 204736 74540
rect 188272 74454 188798 74506
rect 188850 74454 188902 74506
rect 188954 74454 189006 74506
rect 189058 74454 204736 74506
rect 188272 74420 204736 74454
rect 1344 73722 17920 73756
rect 1344 73670 5138 73722
rect 5190 73670 5242 73722
rect 5294 73670 5346 73722
rect 5398 73670 17920 73722
rect 1344 73636 17920 73670
rect 188272 73722 204736 73756
rect 188272 73670 189458 73722
rect 189510 73670 189562 73722
rect 189614 73670 189666 73722
rect 189718 73670 204736 73722
rect 188272 73636 204736 73670
rect 17502 73218 17554 73230
rect 17502 73154 17554 73166
rect 1344 72938 17920 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 17920 72938
rect 1344 72852 17920 72886
rect 188272 72938 204736 72972
rect 188272 72886 188798 72938
rect 188850 72886 188902 72938
rect 188954 72886 189006 72938
rect 189058 72886 204736 72938
rect 188272 72852 204736 72886
rect 1344 72154 17920 72188
rect 1344 72102 5138 72154
rect 5190 72102 5242 72154
rect 5294 72102 5346 72154
rect 5398 72102 17920 72154
rect 1344 72068 17920 72102
rect 188272 72154 204736 72188
rect 188272 72102 189458 72154
rect 189510 72102 189562 72154
rect 189614 72102 189666 72154
rect 189718 72102 204736 72154
rect 188272 72068 204736 72102
rect 1344 71370 17920 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 17920 71370
rect 1344 71284 17920 71318
rect 188272 71370 204736 71404
rect 188272 71318 188798 71370
rect 188850 71318 188902 71370
rect 188954 71318 189006 71370
rect 189058 71318 204736 71370
rect 188272 71284 204736 71318
rect 1710 71090 1762 71102
rect 1710 71026 1762 71038
rect 1344 70586 17920 70620
rect 1344 70534 5138 70586
rect 5190 70534 5242 70586
rect 5294 70534 5346 70586
rect 5398 70534 17920 70586
rect 1344 70500 17920 70534
rect 188272 70586 204736 70620
rect 188272 70534 189458 70586
rect 189510 70534 189562 70586
rect 189614 70534 189666 70586
rect 189718 70534 204736 70586
rect 188272 70500 204736 70534
rect 1344 69802 17920 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 17920 69802
rect 1344 69716 17920 69750
rect 188272 69802 204736 69836
rect 188272 69750 188798 69802
rect 188850 69750 188902 69802
rect 188954 69750 189006 69802
rect 189058 69750 204736 69802
rect 188272 69716 204736 69750
rect 1344 69018 17920 69052
rect 1344 68966 5138 69018
rect 5190 68966 5242 69018
rect 5294 68966 5346 69018
rect 5398 68966 17920 69018
rect 1344 68932 17920 68966
rect 188272 69018 204736 69052
rect 188272 68966 189458 69018
rect 189510 68966 189562 69018
rect 189614 68966 189666 69018
rect 189718 68966 204736 69018
rect 188272 68932 204736 68966
rect 1344 68234 17920 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 17920 68234
rect 1344 68148 17920 68182
rect 188272 68234 204736 68268
rect 188272 68182 188798 68234
rect 188850 68182 188902 68234
rect 188954 68182 189006 68234
rect 189058 68182 204736 68234
rect 188272 68148 204736 68182
rect 1344 67450 17920 67484
rect 1344 67398 5138 67450
rect 5190 67398 5242 67450
rect 5294 67398 5346 67450
rect 5398 67398 17920 67450
rect 1344 67364 17920 67398
rect 188272 67450 204736 67484
rect 188272 67398 189458 67450
rect 189510 67398 189562 67450
rect 189614 67398 189666 67450
rect 189718 67398 204736 67450
rect 188272 67364 204736 67398
rect 2034 67118 2046 67170
rect 2098 67118 2110 67170
rect 1710 67058 1762 67070
rect 201170 67006 201182 67058
rect 201234 67006 201246 67058
rect 1710 66994 1762 67006
rect 2494 66946 2546 66958
rect 203186 66894 203198 66946
rect 203250 66894 203262 66946
rect 2494 66882 2546 66894
rect 1344 66666 17920 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 17920 66666
rect 1344 66580 17920 66614
rect 188272 66666 204736 66700
rect 188272 66614 188798 66666
rect 188850 66614 188902 66666
rect 188954 66614 189006 66666
rect 189058 66614 204736 66666
rect 188272 66580 204736 66614
rect 203982 66386 204034 66398
rect 203982 66322 204034 66334
rect 1344 65882 17920 65916
rect 1344 65830 5138 65882
rect 5190 65830 5242 65882
rect 5294 65830 5346 65882
rect 5398 65830 17920 65882
rect 1344 65796 17920 65830
rect 188272 65882 204736 65916
rect 188272 65830 189458 65882
rect 189510 65830 189562 65882
rect 189614 65830 189666 65882
rect 189718 65830 204736 65882
rect 188272 65796 204736 65830
rect 1344 65098 17920 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 17920 65098
rect 1344 65012 17920 65046
rect 188272 65098 204736 65132
rect 188272 65046 188798 65098
rect 188850 65046 188902 65098
rect 188954 65046 189006 65098
rect 189058 65046 204736 65098
rect 188272 65012 204736 65046
rect 1344 64314 17920 64348
rect 1344 64262 5138 64314
rect 5190 64262 5242 64314
rect 5294 64262 5346 64314
rect 5398 64262 17920 64314
rect 1344 64228 17920 64262
rect 188272 64314 204736 64348
rect 188272 64262 189458 64314
rect 189510 64262 189562 64314
rect 189614 64262 189666 64314
rect 189718 64262 204736 64314
rect 188272 64228 204736 64262
rect 1344 63530 17920 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 17920 63530
rect 1344 63444 17920 63478
rect 188272 63530 204736 63564
rect 188272 63478 188798 63530
rect 188850 63478 188902 63530
rect 188954 63478 189006 63530
rect 189058 63478 204736 63530
rect 188272 63444 204736 63478
rect 1710 62914 1762 62926
rect 1710 62850 1762 62862
rect 1344 62746 17920 62780
rect 1344 62694 5138 62746
rect 5190 62694 5242 62746
rect 5294 62694 5346 62746
rect 5398 62694 17920 62746
rect 1344 62660 17920 62694
rect 188272 62746 204736 62780
rect 188272 62694 189458 62746
rect 189510 62694 189562 62746
rect 189614 62694 189666 62746
rect 189718 62694 204736 62746
rect 188272 62660 204736 62694
rect 1344 61962 17920 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 17920 61962
rect 1344 61876 17920 61910
rect 188272 61962 204736 61996
rect 188272 61910 188798 61962
rect 188850 61910 188902 61962
rect 188954 61910 189006 61962
rect 189058 61910 204736 61962
rect 188272 61876 204736 61910
rect 1344 61178 17920 61212
rect 1344 61126 5138 61178
rect 5190 61126 5242 61178
rect 5294 61126 5346 61178
rect 5398 61126 17920 61178
rect 1344 61092 17920 61126
rect 188272 61178 204736 61212
rect 188272 61126 189458 61178
rect 189510 61126 189562 61178
rect 189614 61126 189666 61178
rect 189718 61126 204736 61178
rect 188272 61092 204736 61126
rect 1344 60394 17920 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 17920 60394
rect 1344 60308 17920 60342
rect 188272 60394 204736 60428
rect 188272 60342 188798 60394
rect 188850 60342 188902 60394
rect 188954 60342 189006 60394
rect 189058 60342 204736 60394
rect 188272 60308 204736 60342
rect 1344 59610 17920 59644
rect 1344 59558 5138 59610
rect 5190 59558 5242 59610
rect 5294 59558 5346 59610
rect 5398 59558 17920 59610
rect 1344 59524 17920 59558
rect 188272 59610 204736 59644
rect 188272 59558 189458 59610
rect 189510 59558 189562 59610
rect 189614 59558 189666 59610
rect 189718 59558 204736 59610
rect 188272 59524 204736 59558
rect 1710 58994 1762 59006
rect 1710 58930 1762 58942
rect 1344 58826 17920 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 17920 58826
rect 1344 58740 17920 58774
rect 188272 58826 204736 58860
rect 188272 58774 188798 58826
rect 188850 58774 188902 58826
rect 188954 58774 189006 58826
rect 189058 58774 204736 58826
rect 188272 58740 204736 58774
rect 1344 58042 17920 58076
rect 1344 57990 5138 58042
rect 5190 57990 5242 58042
rect 5294 57990 5346 58042
rect 5398 57990 17920 58042
rect 1344 57956 17920 57990
rect 188272 58042 204736 58076
rect 188272 57990 189458 58042
rect 189510 57990 189562 58042
rect 189614 57990 189666 58042
rect 189718 57990 204736 58042
rect 188272 57956 204736 57990
rect 1344 57258 17920 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 17920 57258
rect 1344 57172 17920 57206
rect 188272 57258 204736 57292
rect 188272 57206 188798 57258
rect 188850 57206 188902 57258
rect 188954 57206 189006 57258
rect 189058 57206 204736 57258
rect 188272 57172 204736 57206
rect 1344 56474 17920 56508
rect 1344 56422 5138 56474
rect 5190 56422 5242 56474
rect 5294 56422 5346 56474
rect 5398 56422 17920 56474
rect 1344 56388 17920 56422
rect 188272 56474 204736 56508
rect 188272 56422 189458 56474
rect 189510 56422 189562 56474
rect 189614 56422 189666 56474
rect 189718 56422 204736 56474
rect 188272 56388 204736 56422
rect 1344 55690 17920 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 17920 55690
rect 1344 55604 17920 55638
rect 188272 55690 204736 55724
rect 188272 55638 188798 55690
rect 188850 55638 188902 55690
rect 188954 55638 189006 55690
rect 189058 55638 204736 55690
rect 188272 55604 204736 55638
rect 2270 55298 2322 55310
rect 2270 55234 2322 55246
rect 1710 55186 1762 55198
rect 1710 55122 1762 55134
rect 1344 54906 17920 54940
rect 1344 54854 5138 54906
rect 5190 54854 5242 54906
rect 5294 54854 5346 54906
rect 5398 54854 17920 54906
rect 1344 54820 17920 54854
rect 188272 54906 204736 54940
rect 188272 54854 189458 54906
rect 189510 54854 189562 54906
rect 189614 54854 189666 54906
rect 189718 54854 204736 54906
rect 188272 54820 204736 54854
rect 1822 54738 1874 54750
rect 1822 54674 1874 54686
rect 1344 54122 17920 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 17920 54122
rect 1344 54036 17920 54070
rect 188272 54122 204736 54156
rect 188272 54070 188798 54122
rect 188850 54070 188902 54122
rect 188954 54070 189006 54122
rect 189058 54070 204736 54122
rect 188272 54036 204736 54070
rect 1344 53338 17920 53372
rect 1344 53286 5138 53338
rect 5190 53286 5242 53338
rect 5294 53286 5346 53338
rect 5398 53286 17920 53338
rect 1344 53252 17920 53286
rect 188272 53338 204736 53372
rect 188272 53286 189458 53338
rect 189510 53286 189562 53338
rect 189614 53286 189666 53338
rect 189718 53286 204736 53338
rect 188272 53252 204736 53286
rect 1344 52554 17920 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 17920 52554
rect 1344 52468 17920 52502
rect 188272 52554 204736 52588
rect 188272 52502 188798 52554
rect 188850 52502 188902 52554
rect 188954 52502 189006 52554
rect 189058 52502 204736 52554
rect 188272 52468 204736 52502
rect 1710 51938 1762 51950
rect 1710 51874 1762 51886
rect 1344 51770 17920 51804
rect 1344 51718 5138 51770
rect 5190 51718 5242 51770
rect 5294 51718 5346 51770
rect 5398 51718 17920 51770
rect 1344 51684 17920 51718
rect 188272 51770 204736 51804
rect 188272 51718 189458 51770
rect 189510 51718 189562 51770
rect 189614 51718 189666 51770
rect 189718 51718 204736 51770
rect 188272 51684 204736 51718
rect 1344 50986 17920 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 17920 50986
rect 1344 50900 17920 50934
rect 188272 50986 204736 51020
rect 188272 50934 188798 50986
rect 188850 50934 188902 50986
rect 188954 50934 189006 50986
rect 189058 50934 204736 50986
rect 188272 50900 204736 50934
rect 1344 50202 17920 50236
rect 1344 50150 5138 50202
rect 5190 50150 5242 50202
rect 5294 50150 5346 50202
rect 5398 50150 17920 50202
rect 1344 50116 17920 50150
rect 188272 50202 204736 50236
rect 188272 50150 189458 50202
rect 189510 50150 189562 50202
rect 189614 50150 189666 50202
rect 189718 50150 204736 50202
rect 188272 50116 204736 50150
rect 203758 49922 203810 49934
rect 203758 49858 203810 49870
rect 1344 49418 17920 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 17920 49418
rect 1344 49332 17920 49366
rect 188272 49418 204736 49452
rect 188272 49366 188798 49418
rect 188850 49366 188902 49418
rect 188954 49366 189006 49418
rect 189058 49366 204736 49418
rect 188272 49332 204736 49366
rect 1344 48634 17920 48668
rect 1344 48582 5138 48634
rect 5190 48582 5242 48634
rect 5294 48582 5346 48634
rect 5398 48582 17920 48634
rect 1344 48548 17920 48582
rect 188272 48634 204736 48668
rect 188272 48582 189458 48634
rect 189510 48582 189562 48634
rect 189614 48582 189666 48634
rect 189718 48582 204736 48634
rect 188272 48548 204736 48582
rect 1710 48018 1762 48030
rect 1710 47954 1762 47966
rect 1344 47850 17920 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 17920 47850
rect 1344 47764 17920 47798
rect 188272 47850 204736 47884
rect 188272 47798 188798 47850
rect 188850 47798 188902 47850
rect 188954 47798 189006 47850
rect 189058 47798 204736 47850
rect 188272 47764 204736 47798
rect 173954 47182 173966 47234
rect 174018 47231 174030 47234
rect 174402 47231 174414 47234
rect 174018 47185 174414 47231
rect 174018 47182 174030 47185
rect 174402 47182 174414 47185
rect 174466 47182 174478 47234
rect 1344 47066 17920 47100
rect 1344 47014 5138 47066
rect 5190 47014 5242 47066
rect 5294 47014 5346 47066
rect 5398 47014 17920 47066
rect 1344 46980 17920 47014
rect 188272 47066 204736 47100
rect 188272 47014 189458 47066
rect 189510 47014 189562 47066
rect 189614 47014 189666 47066
rect 189718 47014 204736 47066
rect 188272 46980 204736 47014
rect 1344 46282 17920 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 17920 46282
rect 1344 46196 17920 46230
rect 188272 46282 204736 46316
rect 188272 46230 188798 46282
rect 188850 46230 188902 46282
rect 188954 46230 189006 46282
rect 189058 46230 204736 46282
rect 188272 46196 204736 46230
rect 1344 45498 17920 45532
rect 1344 45446 5138 45498
rect 5190 45446 5242 45498
rect 5294 45446 5346 45498
rect 5398 45446 17920 45498
rect 1344 45412 17920 45446
rect 188272 45498 204736 45532
rect 188272 45446 189458 45498
rect 189510 45446 189562 45498
rect 189614 45446 189666 45498
rect 189718 45446 204736 45498
rect 188272 45412 204736 45446
rect 1344 44714 17920 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 17920 44714
rect 1344 44628 17920 44662
rect 188272 44714 204736 44748
rect 188272 44662 188798 44714
rect 188850 44662 188902 44714
rect 188954 44662 189006 44714
rect 189058 44662 204736 44714
rect 188272 44628 204736 44662
rect 2270 44322 2322 44334
rect 1810 44270 1822 44322
rect 1874 44270 1886 44322
rect 2270 44258 2322 44270
rect 1344 43930 17920 43964
rect 1344 43878 5138 43930
rect 5190 43878 5242 43930
rect 5294 43878 5346 43930
rect 5398 43878 17920 43930
rect 1344 43844 17920 43878
rect 188272 43930 204736 43964
rect 188272 43878 189458 43930
rect 189510 43878 189562 43930
rect 189614 43878 189666 43930
rect 189718 43878 204736 43930
rect 188272 43844 204736 43878
rect 1822 43762 1874 43774
rect 1822 43698 1874 43710
rect 1344 43146 17920 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 17920 43146
rect 1344 43060 17920 43094
rect 188272 43146 204736 43180
rect 188272 43094 188798 43146
rect 188850 43094 188902 43146
rect 188954 43094 189006 43146
rect 189058 43094 204736 43146
rect 188272 43060 204736 43094
rect 1344 42362 17920 42396
rect 1344 42310 5138 42362
rect 5190 42310 5242 42362
rect 5294 42310 5346 42362
rect 5398 42310 17920 42362
rect 1344 42276 17920 42310
rect 188272 42362 204736 42396
rect 188272 42310 189458 42362
rect 189510 42310 189562 42362
rect 189614 42310 189666 42362
rect 189718 42310 204736 42362
rect 188272 42276 204736 42310
rect 1344 41578 17920 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 17920 41578
rect 1344 41492 17920 41526
rect 188272 41578 204736 41612
rect 188272 41526 188798 41578
rect 188850 41526 188902 41578
rect 188954 41526 189006 41578
rect 189058 41526 204736 41578
rect 188272 41492 204736 41526
rect 204094 41298 204146 41310
rect 204094 41234 204146 41246
rect 201730 41134 201742 41186
rect 201794 41134 201806 41186
rect 201406 40962 201458 40974
rect 201406 40898 201458 40910
rect 1344 40794 17920 40828
rect 1344 40742 5138 40794
rect 5190 40742 5242 40794
rect 5294 40742 5346 40794
rect 5398 40742 17920 40794
rect 1344 40708 17920 40742
rect 188272 40794 204736 40828
rect 188272 40742 189458 40794
rect 189510 40742 189562 40794
rect 189614 40742 189666 40794
rect 189718 40742 204736 40794
rect 188272 40708 204736 40742
rect 1710 40514 1762 40526
rect 1710 40450 1762 40462
rect 1344 40010 17920 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 17920 40010
rect 1344 39924 17920 39958
rect 188272 40010 204736 40044
rect 188272 39958 188798 40010
rect 188850 39958 188902 40010
rect 188954 39958 189006 40010
rect 189058 39958 204736 40010
rect 188272 39924 204736 39958
rect 1344 39226 17920 39260
rect 1344 39174 5138 39226
rect 5190 39174 5242 39226
rect 5294 39174 5346 39226
rect 5398 39174 17920 39226
rect 1344 39140 17920 39174
rect 188272 39226 204736 39260
rect 188272 39174 189458 39226
rect 189510 39174 189562 39226
rect 189614 39174 189666 39226
rect 189718 39174 204736 39226
rect 188272 39140 204736 39174
rect 188750 38722 188802 38734
rect 188750 38658 188802 38670
rect 1344 38442 17920 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 17920 38442
rect 1344 38356 17920 38390
rect 188272 38442 204736 38476
rect 188272 38390 188798 38442
rect 188850 38390 188902 38442
rect 188954 38390 189006 38442
rect 189058 38390 204736 38442
rect 188272 38356 204736 38390
rect 1344 37658 17920 37692
rect 1344 37606 5138 37658
rect 5190 37606 5242 37658
rect 5294 37606 5346 37658
rect 5398 37606 17920 37658
rect 1344 37572 17920 37606
rect 188272 37658 204736 37692
rect 188272 37606 189458 37658
rect 189510 37606 189562 37658
rect 189614 37606 189666 37658
rect 189718 37606 204736 37658
rect 188272 37572 204736 37606
rect 1344 36874 17920 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 17920 36874
rect 1344 36788 17920 36822
rect 188272 36874 204736 36908
rect 188272 36822 188798 36874
rect 188850 36822 188902 36874
rect 188954 36822 189006 36874
rect 189058 36822 204736 36874
rect 188272 36788 204736 36822
rect 1710 36594 1762 36606
rect 1710 36530 1762 36542
rect 17614 36258 17666 36270
rect 17614 36194 17666 36206
rect 1344 36090 17920 36124
rect 1344 36038 5138 36090
rect 5190 36038 5242 36090
rect 5294 36038 5346 36090
rect 5398 36038 17920 36090
rect 1344 36004 17920 36038
rect 188272 36090 204736 36124
rect 188272 36038 189458 36090
rect 189510 36038 189562 36090
rect 189614 36038 189666 36090
rect 189718 36038 204736 36090
rect 188272 36004 204736 36038
rect 16942 35586 16994 35598
rect 16942 35522 16994 35534
rect 17614 35586 17666 35598
rect 17614 35522 17666 35534
rect 1344 35306 17920 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 17920 35306
rect 1344 35220 17920 35254
rect 188272 35306 204736 35340
rect 188272 35254 188798 35306
rect 188850 35254 188902 35306
rect 188954 35254 189006 35306
rect 189058 35254 204736 35306
rect 188272 35220 204736 35254
rect 1344 34522 17920 34556
rect 1344 34470 5138 34522
rect 5190 34470 5242 34522
rect 5294 34470 5346 34522
rect 5398 34470 17920 34522
rect 1344 34436 17920 34470
rect 188272 34522 204736 34556
rect 188272 34470 189458 34522
rect 189510 34470 189562 34522
rect 189614 34470 189666 34522
rect 189718 34470 204736 34522
rect 188272 34436 204736 34470
rect 1344 33738 17920 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 17920 33738
rect 1344 33652 17920 33686
rect 188272 33738 204736 33772
rect 188272 33686 188798 33738
rect 188850 33686 188902 33738
rect 188954 33686 189006 33738
rect 189058 33686 204736 33738
rect 188272 33652 204736 33686
rect 1344 32954 17920 32988
rect 1344 32902 5138 32954
rect 5190 32902 5242 32954
rect 5294 32902 5346 32954
rect 5398 32902 17920 32954
rect 1344 32868 17920 32902
rect 188272 32954 204736 32988
rect 188272 32902 189458 32954
rect 189510 32902 189562 32954
rect 189614 32902 189666 32954
rect 189718 32902 204736 32954
rect 188272 32868 204736 32902
rect 2046 32786 2098 32798
rect 2046 32722 2098 32734
rect 1710 32562 1762 32574
rect 1710 32498 1762 32510
rect 2494 32450 2546 32462
rect 2494 32386 2546 32398
rect 1344 32170 17920 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 17920 32170
rect 1344 32084 17920 32118
rect 188272 32170 204736 32204
rect 188272 32118 188798 32170
rect 188850 32118 188902 32170
rect 188954 32118 189006 32170
rect 189058 32118 204736 32170
rect 188272 32084 204736 32118
rect 1344 31386 17920 31420
rect 1344 31334 5138 31386
rect 5190 31334 5242 31386
rect 5294 31334 5346 31386
rect 5398 31334 17920 31386
rect 1344 31300 17920 31334
rect 188272 31386 204736 31420
rect 188272 31334 189458 31386
rect 189510 31334 189562 31386
rect 189614 31334 189666 31386
rect 189718 31334 204736 31386
rect 188272 31300 204736 31334
rect 1344 30602 17920 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 17920 30602
rect 1344 30516 17920 30550
rect 188272 30602 204736 30636
rect 188272 30550 188798 30602
rect 188850 30550 188902 30602
rect 188954 30550 189006 30602
rect 189058 30550 204736 30602
rect 188272 30516 204736 30550
rect 1344 29818 17920 29852
rect 1344 29766 5138 29818
rect 5190 29766 5242 29818
rect 5294 29766 5346 29818
rect 5398 29766 17920 29818
rect 1344 29732 17920 29766
rect 188272 29818 204736 29852
rect 188272 29766 189458 29818
rect 189510 29766 189562 29818
rect 189614 29766 189666 29818
rect 189718 29766 204736 29818
rect 188272 29732 204736 29766
rect 1344 29034 17920 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 17920 29034
rect 1344 28948 17920 28982
rect 188272 29034 204736 29068
rect 188272 28982 188798 29034
rect 188850 28982 188902 29034
rect 188954 28982 189006 29034
rect 189058 28982 204736 29034
rect 188272 28948 204736 28982
rect 1710 28530 1762 28542
rect 1710 28466 1762 28478
rect 1344 28250 17920 28284
rect 1344 28198 5138 28250
rect 5190 28198 5242 28250
rect 5294 28198 5346 28250
rect 5398 28198 17920 28250
rect 1344 28164 17920 28198
rect 188272 28250 204736 28284
rect 188272 28198 189458 28250
rect 189510 28198 189562 28250
rect 189614 28198 189666 28250
rect 189718 28198 204736 28250
rect 188272 28164 204736 28198
rect 1344 27466 17920 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 17920 27466
rect 1344 27380 17920 27414
rect 188272 27466 204736 27500
rect 188272 27414 188798 27466
rect 188850 27414 188902 27466
rect 188954 27414 189006 27466
rect 189058 27414 204736 27466
rect 188272 27380 204736 27414
rect 1344 26682 17920 26716
rect 1344 26630 5138 26682
rect 5190 26630 5242 26682
rect 5294 26630 5346 26682
rect 5398 26630 17920 26682
rect 1344 26596 17920 26630
rect 188272 26682 204736 26716
rect 188272 26630 189458 26682
rect 189510 26630 189562 26682
rect 189614 26630 189666 26682
rect 189718 26630 204736 26682
rect 188272 26596 204736 26630
rect 1344 25898 17920 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 17920 25898
rect 1344 25812 17920 25846
rect 188272 25898 204736 25932
rect 188272 25846 188798 25898
rect 188850 25846 188902 25898
rect 188954 25846 189006 25898
rect 189058 25846 204736 25898
rect 188272 25812 204736 25846
rect 1710 25618 1762 25630
rect 1710 25554 1762 25566
rect 1344 25114 17920 25148
rect 1344 25062 5138 25114
rect 5190 25062 5242 25114
rect 5294 25062 5346 25114
rect 5398 25062 17920 25114
rect 1344 25028 17920 25062
rect 188272 25114 204736 25148
rect 188272 25062 189458 25114
rect 189510 25062 189562 25114
rect 189614 25062 189666 25114
rect 189718 25062 204736 25114
rect 188272 25028 204736 25062
rect 1344 24330 17920 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 17920 24330
rect 1344 24244 17920 24278
rect 188272 24330 204736 24364
rect 188272 24278 188798 24330
rect 188850 24278 188902 24330
rect 188954 24278 189006 24330
rect 189058 24278 204736 24330
rect 188272 24244 204736 24278
rect 204318 23714 204370 23726
rect 204318 23650 204370 23662
rect 1344 23546 17920 23580
rect 1344 23494 5138 23546
rect 5190 23494 5242 23546
rect 5294 23494 5346 23546
rect 5398 23494 17920 23546
rect 1344 23460 17920 23494
rect 188272 23546 204736 23580
rect 188272 23494 189458 23546
rect 189510 23494 189562 23546
rect 189614 23494 189666 23546
rect 189718 23494 204736 23546
rect 188272 23460 204736 23494
rect 1344 22762 17920 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 17920 22762
rect 1344 22676 17920 22710
rect 188272 22762 204736 22796
rect 188272 22710 188798 22762
rect 188850 22710 188902 22762
rect 188954 22710 189006 22762
rect 189058 22710 204736 22762
rect 188272 22676 204736 22710
rect 1344 21978 17920 22012
rect 1344 21926 5138 21978
rect 5190 21926 5242 21978
rect 5294 21926 5346 21978
rect 5398 21926 17920 21978
rect 1344 21892 17920 21926
rect 188272 21978 204736 22012
rect 188272 21926 189458 21978
rect 189510 21926 189562 21978
rect 189614 21926 189666 21978
rect 189718 21926 204736 21978
rect 188272 21892 204736 21926
rect 2046 21810 2098 21822
rect 2046 21746 2098 21758
rect 1710 21586 1762 21598
rect 1710 21522 1762 21534
rect 2494 21474 2546 21486
rect 2494 21410 2546 21422
rect 1344 21194 17920 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 17920 21194
rect 1344 21108 17920 21142
rect 188272 21194 204736 21228
rect 188272 21142 188798 21194
rect 188850 21142 188902 21194
rect 188954 21142 189006 21194
rect 189058 21142 204736 21194
rect 188272 21108 204736 21142
rect 1344 20410 17920 20444
rect 1344 20358 5138 20410
rect 5190 20358 5242 20410
rect 5294 20358 5346 20410
rect 5398 20358 17920 20410
rect 1344 20324 17920 20358
rect 188272 20410 204736 20444
rect 188272 20358 189458 20410
rect 189510 20358 189562 20410
rect 189614 20358 189666 20410
rect 189718 20358 204736 20410
rect 188272 20324 204736 20358
rect 1344 19626 17920 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 17920 19626
rect 1344 19540 17920 19574
rect 188272 19626 204736 19660
rect 188272 19574 188798 19626
rect 188850 19574 188902 19626
rect 188954 19574 189006 19626
rect 189058 19574 204736 19626
rect 188272 19540 204736 19574
rect 1344 18842 17920 18876
rect 1344 18790 5138 18842
rect 5190 18790 5242 18842
rect 5294 18790 5346 18842
rect 5398 18790 17920 18842
rect 1344 18756 17920 18790
rect 188272 18842 204736 18876
rect 188272 18790 189458 18842
rect 189510 18790 189562 18842
rect 189614 18790 189666 18842
rect 189718 18790 204736 18842
rect 188272 18756 204736 18790
rect 1344 18058 17920 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 17920 18058
rect 1344 17972 17920 18006
rect 188272 18058 204736 18092
rect 188272 18006 188798 18058
rect 188850 18006 188902 18058
rect 188954 18006 189006 18058
rect 189058 18006 204736 18058
rect 188272 17972 204736 18006
rect 1710 17442 1762 17454
rect 1710 17378 1762 17390
rect 1344 17274 204736 17308
rect 1344 17222 5138 17274
rect 5190 17222 5242 17274
rect 5294 17222 5346 17274
rect 5398 17222 35858 17274
rect 35910 17222 35962 17274
rect 36014 17222 36066 17274
rect 36118 17222 66578 17274
rect 66630 17222 66682 17274
rect 66734 17222 66786 17274
rect 66838 17222 97298 17274
rect 97350 17222 97402 17274
rect 97454 17222 97506 17274
rect 97558 17222 128018 17274
rect 128070 17222 128122 17274
rect 128174 17222 128226 17274
rect 128278 17222 158738 17274
rect 158790 17222 158842 17274
rect 158894 17222 158946 17274
rect 158998 17222 189458 17274
rect 189510 17222 189562 17274
rect 189614 17222 189666 17274
rect 189718 17222 204736 17274
rect 1344 17188 204736 17222
rect 44718 17106 44770 17118
rect 44718 17042 44770 17054
rect 48190 17106 48242 17118
rect 48190 17042 48242 17054
rect 51550 17106 51602 17118
rect 51550 17042 51602 17054
rect 55134 17106 55186 17118
rect 55134 17042 55186 17054
rect 59054 17106 59106 17118
rect 59054 17042 59106 17054
rect 61966 17106 62018 17118
rect 61966 17042 62018 17054
rect 65438 17106 65490 17118
rect 65438 17042 65490 17054
rect 68798 17106 68850 17118
rect 68798 17042 68850 17054
rect 72158 17106 72210 17118
rect 72158 17042 72210 17054
rect 75518 17106 75570 17118
rect 75518 17042 75570 17054
rect 78990 17106 79042 17118
rect 78990 17042 79042 17054
rect 82350 17106 82402 17118
rect 82350 17042 82402 17054
rect 82910 17106 82962 17118
rect 82910 17042 82962 17054
rect 97134 17106 97186 17118
rect 97134 17042 97186 17054
rect 111246 17106 111298 17118
rect 111246 17042 111298 17054
rect 140030 17106 140082 17118
rect 140030 17042 140082 17054
rect 154366 17106 154418 17118
rect 154366 17042 154418 17054
rect 67902 16882 67954 16894
rect 67902 16818 67954 16830
rect 125582 16882 125634 16894
rect 125582 16818 125634 16830
rect 1344 16490 204736 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 127358 16490
rect 127410 16438 127462 16490
rect 127514 16438 127566 16490
rect 127618 16438 158078 16490
rect 158130 16438 158182 16490
rect 158234 16438 158286 16490
rect 158338 16438 188798 16490
rect 188850 16438 188902 16490
rect 188954 16438 189006 16490
rect 189058 16438 204736 16490
rect 1344 16404 204736 16438
rect 1344 15706 204736 15740
rect 1344 15654 5138 15706
rect 5190 15654 5242 15706
rect 5294 15654 5346 15706
rect 5398 15654 35858 15706
rect 35910 15654 35962 15706
rect 36014 15654 36066 15706
rect 36118 15654 66578 15706
rect 66630 15654 66682 15706
rect 66734 15654 66786 15706
rect 66838 15654 97298 15706
rect 97350 15654 97402 15706
rect 97454 15654 97506 15706
rect 97558 15654 128018 15706
rect 128070 15654 128122 15706
rect 128174 15654 128226 15706
rect 128278 15654 158738 15706
rect 158790 15654 158842 15706
rect 158894 15654 158946 15706
rect 158998 15654 189458 15706
rect 189510 15654 189562 15706
rect 189614 15654 189666 15706
rect 189718 15654 204736 15706
rect 1344 15620 204736 15654
rect 1344 14922 204736 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 127358 14922
rect 127410 14870 127462 14922
rect 127514 14870 127566 14922
rect 127618 14870 158078 14922
rect 158130 14870 158182 14922
rect 158234 14870 158286 14922
rect 158338 14870 188798 14922
rect 188850 14870 188902 14922
rect 188954 14870 189006 14922
rect 189058 14870 204736 14922
rect 1344 14836 204736 14870
rect 204094 14642 204146 14654
rect 204094 14578 204146 14590
rect 201730 14478 201742 14530
rect 201794 14478 201806 14530
rect 1344 14138 204736 14172
rect 1344 14086 5138 14138
rect 5190 14086 5242 14138
rect 5294 14086 5346 14138
rect 5398 14086 35858 14138
rect 35910 14086 35962 14138
rect 36014 14086 36066 14138
rect 36118 14086 66578 14138
rect 66630 14086 66682 14138
rect 66734 14086 66786 14138
rect 66838 14086 97298 14138
rect 97350 14086 97402 14138
rect 97454 14086 97506 14138
rect 97558 14086 128018 14138
rect 128070 14086 128122 14138
rect 128174 14086 128226 14138
rect 128278 14086 158738 14138
rect 158790 14086 158842 14138
rect 158894 14086 158946 14138
rect 158998 14086 189458 14138
rect 189510 14086 189562 14138
rect 189614 14086 189666 14138
rect 189718 14086 204736 14138
rect 1344 14052 204736 14086
rect 204318 13970 204370 13982
rect 204318 13906 204370 13918
rect 1710 13522 1762 13534
rect 1710 13458 1762 13470
rect 1344 13354 204736 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 127358 13354
rect 127410 13302 127462 13354
rect 127514 13302 127566 13354
rect 127618 13302 158078 13354
rect 158130 13302 158182 13354
rect 158234 13302 158286 13354
rect 158338 13302 188798 13354
rect 188850 13302 188902 13354
rect 188954 13302 189006 13354
rect 189058 13302 204736 13354
rect 1344 13268 204736 13302
rect 1344 12570 204736 12604
rect 1344 12518 5138 12570
rect 5190 12518 5242 12570
rect 5294 12518 5346 12570
rect 5398 12518 35858 12570
rect 35910 12518 35962 12570
rect 36014 12518 36066 12570
rect 36118 12518 66578 12570
rect 66630 12518 66682 12570
rect 66734 12518 66786 12570
rect 66838 12518 97298 12570
rect 97350 12518 97402 12570
rect 97454 12518 97506 12570
rect 97558 12518 128018 12570
rect 128070 12518 128122 12570
rect 128174 12518 128226 12570
rect 128278 12518 158738 12570
rect 158790 12518 158842 12570
rect 158894 12518 158946 12570
rect 158998 12518 189458 12570
rect 189510 12518 189562 12570
rect 189614 12518 189666 12570
rect 189718 12518 204736 12570
rect 1344 12484 204736 12518
rect 1344 11786 204736 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 127358 11786
rect 127410 11734 127462 11786
rect 127514 11734 127566 11786
rect 127618 11734 158078 11786
rect 158130 11734 158182 11786
rect 158234 11734 158286 11786
rect 158338 11734 188798 11786
rect 188850 11734 188902 11786
rect 188954 11734 189006 11786
rect 189058 11734 204736 11786
rect 1344 11700 204736 11734
rect 1344 11002 204736 11036
rect 1344 10950 5138 11002
rect 5190 10950 5242 11002
rect 5294 10950 5346 11002
rect 5398 10950 35858 11002
rect 35910 10950 35962 11002
rect 36014 10950 36066 11002
rect 36118 10950 66578 11002
rect 66630 10950 66682 11002
rect 66734 10950 66786 11002
rect 66838 10950 97298 11002
rect 97350 10950 97402 11002
rect 97454 10950 97506 11002
rect 97558 10950 128018 11002
rect 128070 10950 128122 11002
rect 128174 10950 128226 11002
rect 128278 10950 158738 11002
rect 158790 10950 158842 11002
rect 158894 10950 158946 11002
rect 158998 10950 189458 11002
rect 189510 10950 189562 11002
rect 189614 10950 189666 11002
rect 189718 10950 204736 11002
rect 1344 10916 204736 10950
rect 1344 10218 204736 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 127358 10218
rect 127410 10166 127462 10218
rect 127514 10166 127566 10218
rect 127618 10166 158078 10218
rect 158130 10166 158182 10218
rect 158234 10166 158286 10218
rect 158338 10166 188798 10218
rect 188850 10166 188902 10218
rect 188954 10166 189006 10218
rect 189058 10166 204736 10218
rect 1344 10132 204736 10166
rect 1710 9602 1762 9614
rect 2494 9602 2546 9614
rect 2034 9550 2046 9602
rect 2098 9550 2110 9602
rect 1710 9538 1762 9550
rect 2494 9538 2546 9550
rect 1344 9434 204736 9468
rect 1344 9382 5138 9434
rect 5190 9382 5242 9434
rect 5294 9382 5346 9434
rect 5398 9382 35858 9434
rect 35910 9382 35962 9434
rect 36014 9382 36066 9434
rect 36118 9382 66578 9434
rect 66630 9382 66682 9434
rect 66734 9382 66786 9434
rect 66838 9382 97298 9434
rect 97350 9382 97402 9434
rect 97454 9382 97506 9434
rect 97558 9382 128018 9434
rect 128070 9382 128122 9434
rect 128174 9382 128226 9434
rect 128278 9382 158738 9434
rect 158790 9382 158842 9434
rect 158894 9382 158946 9434
rect 158998 9382 189458 9434
rect 189510 9382 189562 9434
rect 189614 9382 189666 9434
rect 189718 9382 204736 9434
rect 1344 9348 204736 9382
rect 1344 8650 204736 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 127358 8650
rect 127410 8598 127462 8650
rect 127514 8598 127566 8650
rect 127618 8598 158078 8650
rect 158130 8598 158182 8650
rect 158234 8598 158286 8650
rect 158338 8598 188798 8650
rect 188850 8598 188902 8650
rect 188954 8598 189006 8650
rect 189058 8598 204736 8650
rect 1344 8564 204736 8598
rect 1344 7866 204736 7900
rect 1344 7814 5138 7866
rect 5190 7814 5242 7866
rect 5294 7814 5346 7866
rect 5398 7814 35858 7866
rect 35910 7814 35962 7866
rect 36014 7814 36066 7866
rect 36118 7814 66578 7866
rect 66630 7814 66682 7866
rect 66734 7814 66786 7866
rect 66838 7814 97298 7866
rect 97350 7814 97402 7866
rect 97454 7814 97506 7866
rect 97558 7814 128018 7866
rect 128070 7814 128122 7866
rect 128174 7814 128226 7866
rect 128278 7814 158738 7866
rect 158790 7814 158842 7866
rect 158894 7814 158946 7866
rect 158998 7814 189458 7866
rect 189510 7814 189562 7866
rect 189614 7814 189666 7866
rect 189718 7814 204736 7866
rect 1344 7780 204736 7814
rect 1344 7082 204736 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 127358 7082
rect 127410 7030 127462 7082
rect 127514 7030 127566 7082
rect 127618 7030 158078 7082
rect 158130 7030 158182 7082
rect 158234 7030 158286 7082
rect 158338 7030 188798 7082
rect 188850 7030 188902 7082
rect 188954 7030 189006 7082
rect 189058 7030 204736 7082
rect 1344 6996 204736 7030
rect 1344 6298 204736 6332
rect 1344 6246 5138 6298
rect 5190 6246 5242 6298
rect 5294 6246 5346 6298
rect 5398 6246 35858 6298
rect 35910 6246 35962 6298
rect 36014 6246 36066 6298
rect 36118 6246 66578 6298
rect 66630 6246 66682 6298
rect 66734 6246 66786 6298
rect 66838 6246 97298 6298
rect 97350 6246 97402 6298
rect 97454 6246 97506 6298
rect 97558 6246 128018 6298
rect 128070 6246 128122 6298
rect 128174 6246 128226 6298
rect 128278 6246 158738 6298
rect 158790 6246 158842 6298
rect 158894 6246 158946 6298
rect 158998 6246 189458 6298
rect 189510 6246 189562 6298
rect 189614 6246 189666 6298
rect 189718 6246 204736 6298
rect 1344 6212 204736 6246
rect 1710 6018 1762 6030
rect 1710 5954 1762 5966
rect 1344 5514 204736 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 127358 5514
rect 127410 5462 127462 5514
rect 127514 5462 127566 5514
rect 127618 5462 158078 5514
rect 158130 5462 158182 5514
rect 158234 5462 158286 5514
rect 158338 5462 188798 5514
rect 188850 5462 188902 5514
rect 188954 5462 189006 5514
rect 189058 5462 204736 5514
rect 1344 5428 204736 5462
rect 1344 4730 204736 4764
rect 1344 4678 5138 4730
rect 5190 4678 5242 4730
rect 5294 4678 5346 4730
rect 5398 4678 35858 4730
rect 35910 4678 35962 4730
rect 36014 4678 36066 4730
rect 36118 4678 66578 4730
rect 66630 4678 66682 4730
rect 66734 4678 66786 4730
rect 66838 4678 97298 4730
rect 97350 4678 97402 4730
rect 97454 4678 97506 4730
rect 97558 4678 128018 4730
rect 128070 4678 128122 4730
rect 128174 4678 128226 4730
rect 128278 4678 158738 4730
rect 158790 4678 158842 4730
rect 158894 4678 158946 4730
rect 158998 4678 189458 4730
rect 189510 4678 189562 4730
rect 189614 4678 189666 4730
rect 189718 4678 204736 4730
rect 1344 4644 204736 4678
rect 1344 3946 204736 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 127358 3946
rect 127410 3894 127462 3946
rect 127514 3894 127566 3946
rect 127618 3894 158078 3946
rect 158130 3894 158182 3946
rect 158234 3894 158286 3946
rect 158338 3894 188798 3946
rect 188850 3894 188902 3946
rect 188954 3894 189006 3946
rect 189058 3894 204736 3946
rect 1344 3860 204736 3894
rect 1710 3666 1762 3678
rect 1710 3602 1762 3614
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 103070 3330 103122 3342
rect 103070 3266 103122 3278
rect 171614 3330 171666 3342
rect 171614 3266 171666 3278
rect 1344 3162 204736 3196
rect 1344 3110 5138 3162
rect 5190 3110 5242 3162
rect 5294 3110 5346 3162
rect 5398 3110 35858 3162
rect 35910 3110 35962 3162
rect 36014 3110 36066 3162
rect 36118 3110 66578 3162
rect 66630 3110 66682 3162
rect 66734 3110 66786 3162
rect 66838 3110 97298 3162
rect 97350 3110 97402 3162
rect 97454 3110 97506 3162
rect 97558 3110 128018 3162
rect 128070 3110 128122 3162
rect 128174 3110 128226 3162
rect 128278 3110 158738 3162
rect 158790 3110 158842 3162
rect 158894 3110 158946 3162
rect 158998 3110 189458 3162
rect 189510 3110 189562 3162
rect 189614 3110 189666 3162
rect 189718 3110 204736 3162
rect 1344 3076 204736 3110
<< via1 >>
rect 133310 157390 133362 157442
rect 134206 157390 134258 157442
rect 87614 157054 87666 157106
rect 88510 157054 88562 157106
rect 89406 157054 89458 157106
rect 156270 157054 156322 157106
rect 157054 157054 157106 157106
rect 157950 157054 158002 157106
rect 5138 156774 5190 156826
rect 5242 156774 5294 156826
rect 5346 156774 5398 156826
rect 35858 156774 35910 156826
rect 35962 156774 36014 156826
rect 36066 156774 36118 156826
rect 66578 156774 66630 156826
rect 66682 156774 66734 156826
rect 66786 156774 66838 156826
rect 97298 156774 97350 156826
rect 97402 156774 97454 156826
rect 97506 156774 97558 156826
rect 128018 156774 128070 156826
rect 128122 156774 128174 156826
rect 128226 156774 128278 156826
rect 158738 156774 158790 156826
rect 158842 156774 158894 156826
rect 158946 156774 158998 156826
rect 189458 156774 189510 156826
rect 189562 156774 189614 156826
rect 189666 156774 189718 156826
rect 11678 156606 11730 156658
rect 19070 156606 19122 156658
rect 19294 156606 19346 156658
rect 34526 156606 34578 156658
rect 43710 156606 43762 156658
rect 57374 156606 57426 156658
rect 66558 156606 66610 156658
rect 80222 156606 80274 156658
rect 89406 156606 89458 156658
rect 103070 156606 103122 156658
rect 110462 156606 110514 156658
rect 110686 156606 110738 156658
rect 125918 156606 125970 156658
rect 135102 156606 135154 156658
rect 148766 156606 148818 156658
rect 157950 156606 158002 156658
rect 163998 156606 164050 156658
rect 186846 156606 186898 156658
rect 1710 156494 1762 156546
rect 87614 156494 87666 156546
rect 41918 156382 41970 156434
rect 64766 156382 64818 156434
rect 88510 156382 88562 156434
rect 134206 156382 134258 156434
rect 157054 156382 157106 156434
rect 2382 156270 2434 156322
rect 20078 156270 20130 156322
rect 42814 156270 42866 156322
rect 65326 156270 65378 156322
rect 111134 156270 111186 156322
rect 156382 156270 156434 156322
rect 4062 156158 4114 156210
rect 26910 156158 26962 156210
rect 49758 156158 49810 156210
rect 72606 156158 72658 156210
rect 95454 156158 95506 156210
rect 118302 156158 118354 156210
rect 133422 156158 133474 156210
rect 141150 156158 141202 156210
rect 4478 155990 4530 156042
rect 4582 155990 4634 156042
rect 4686 155990 4738 156042
rect 35198 155990 35250 156042
rect 35302 155990 35354 156042
rect 35406 155990 35458 156042
rect 65918 155990 65970 156042
rect 66022 155990 66074 156042
rect 66126 155990 66178 156042
rect 96638 155990 96690 156042
rect 96742 155990 96794 156042
rect 96846 155990 96898 156042
rect 127358 155990 127410 156042
rect 127462 155990 127514 156042
rect 127566 155990 127618 156042
rect 158078 155990 158130 156042
rect 158182 155990 158234 156042
rect 158286 155990 158338 156042
rect 188798 155990 188850 156042
rect 188902 155990 188954 156042
rect 189006 155990 189058 156042
rect 171838 155822 171890 155874
rect 1822 155710 1874 155762
rect 194910 155710 194962 155762
rect 174190 155598 174242 155650
rect 196590 155598 196642 155650
rect 174638 155374 174690 155426
rect 197486 155374 197538 155426
rect 5138 155206 5190 155258
rect 5242 155206 5294 155258
rect 5346 155206 5398 155258
rect 35858 155206 35910 155258
rect 35962 155206 36014 155258
rect 36066 155206 36118 155258
rect 66578 155206 66630 155258
rect 66682 155206 66734 155258
rect 66786 155206 66838 155258
rect 97298 155206 97350 155258
rect 97402 155206 97454 155258
rect 97506 155206 97558 155258
rect 128018 155206 128070 155258
rect 128122 155206 128174 155258
rect 128226 155206 128278 155258
rect 158738 155206 158790 155258
rect 158842 155206 158894 155258
rect 158946 155206 158998 155258
rect 189458 155206 189510 155258
rect 189562 155206 189614 155258
rect 189666 155206 189718 155258
rect 1710 154926 1762 154978
rect 204318 154926 204370 154978
rect 4478 154422 4530 154474
rect 4582 154422 4634 154474
rect 4686 154422 4738 154474
rect 35198 154422 35250 154474
rect 35302 154422 35354 154474
rect 35406 154422 35458 154474
rect 65918 154422 65970 154474
rect 66022 154422 66074 154474
rect 66126 154422 66178 154474
rect 96638 154422 96690 154474
rect 96742 154422 96794 154474
rect 96846 154422 96898 154474
rect 127358 154422 127410 154474
rect 127462 154422 127514 154474
rect 127566 154422 127618 154474
rect 158078 154422 158130 154474
rect 158182 154422 158234 154474
rect 158286 154422 158338 154474
rect 188798 154422 188850 154474
rect 188902 154422 188954 154474
rect 189006 154422 189058 154474
rect 5138 153638 5190 153690
rect 5242 153638 5294 153690
rect 5346 153638 5398 153690
rect 35858 153638 35910 153690
rect 35962 153638 36014 153690
rect 36066 153638 36118 153690
rect 66578 153638 66630 153690
rect 66682 153638 66734 153690
rect 66786 153638 66838 153690
rect 97298 153638 97350 153690
rect 97402 153638 97454 153690
rect 97506 153638 97558 153690
rect 128018 153638 128070 153690
rect 128122 153638 128174 153690
rect 128226 153638 128278 153690
rect 158738 153638 158790 153690
rect 158842 153638 158894 153690
rect 158946 153638 158998 153690
rect 189458 153638 189510 153690
rect 189562 153638 189614 153690
rect 189666 153638 189718 153690
rect 4478 152854 4530 152906
rect 4582 152854 4634 152906
rect 4686 152854 4738 152906
rect 35198 152854 35250 152906
rect 35302 152854 35354 152906
rect 35406 152854 35458 152906
rect 65918 152854 65970 152906
rect 66022 152854 66074 152906
rect 66126 152854 66178 152906
rect 96638 152854 96690 152906
rect 96742 152854 96794 152906
rect 96846 152854 96898 152906
rect 127358 152854 127410 152906
rect 127462 152854 127514 152906
rect 127566 152854 127618 152906
rect 158078 152854 158130 152906
rect 158182 152854 158234 152906
rect 158286 152854 158338 152906
rect 188798 152854 188850 152906
rect 188902 152854 188954 152906
rect 189006 152854 189058 152906
rect 5138 152070 5190 152122
rect 5242 152070 5294 152122
rect 5346 152070 5398 152122
rect 35858 152070 35910 152122
rect 35962 152070 36014 152122
rect 36066 152070 36118 152122
rect 66578 152070 66630 152122
rect 66682 152070 66734 152122
rect 66786 152070 66838 152122
rect 97298 152070 97350 152122
rect 97402 152070 97454 152122
rect 97506 152070 97558 152122
rect 128018 152070 128070 152122
rect 128122 152070 128174 152122
rect 128226 152070 128278 152122
rect 158738 152070 158790 152122
rect 158842 152070 158894 152122
rect 158946 152070 158998 152122
rect 189458 152070 189510 152122
rect 189562 152070 189614 152122
rect 189666 152070 189718 152122
rect 4478 151286 4530 151338
rect 4582 151286 4634 151338
rect 4686 151286 4738 151338
rect 35198 151286 35250 151338
rect 35302 151286 35354 151338
rect 35406 151286 35458 151338
rect 65918 151286 65970 151338
rect 66022 151286 66074 151338
rect 66126 151286 66178 151338
rect 96638 151286 96690 151338
rect 96742 151286 96794 151338
rect 96846 151286 96898 151338
rect 127358 151286 127410 151338
rect 127462 151286 127514 151338
rect 127566 151286 127618 151338
rect 158078 151286 158130 151338
rect 158182 151286 158234 151338
rect 158286 151286 158338 151338
rect 188798 151286 188850 151338
rect 188902 151286 188954 151338
rect 189006 151286 189058 151338
rect 1710 151006 1762 151058
rect 5138 150502 5190 150554
rect 5242 150502 5294 150554
rect 5346 150502 5398 150554
rect 35858 150502 35910 150554
rect 35962 150502 36014 150554
rect 36066 150502 36118 150554
rect 66578 150502 66630 150554
rect 66682 150502 66734 150554
rect 66786 150502 66838 150554
rect 97298 150502 97350 150554
rect 97402 150502 97454 150554
rect 97506 150502 97558 150554
rect 128018 150502 128070 150554
rect 128122 150502 128174 150554
rect 128226 150502 128278 150554
rect 158738 150502 158790 150554
rect 158842 150502 158894 150554
rect 158946 150502 158998 150554
rect 189458 150502 189510 150554
rect 189562 150502 189614 150554
rect 189666 150502 189718 150554
rect 4478 149718 4530 149770
rect 4582 149718 4634 149770
rect 4686 149718 4738 149770
rect 35198 149718 35250 149770
rect 35302 149718 35354 149770
rect 35406 149718 35458 149770
rect 65918 149718 65970 149770
rect 66022 149718 66074 149770
rect 66126 149718 66178 149770
rect 96638 149718 96690 149770
rect 96742 149718 96794 149770
rect 96846 149718 96898 149770
rect 127358 149718 127410 149770
rect 127462 149718 127514 149770
rect 127566 149718 127618 149770
rect 158078 149718 158130 149770
rect 158182 149718 158234 149770
rect 158286 149718 158338 149770
rect 188798 149718 188850 149770
rect 188902 149718 188954 149770
rect 189006 149718 189058 149770
rect 5138 148934 5190 148986
rect 5242 148934 5294 148986
rect 5346 148934 5398 148986
rect 35858 148934 35910 148986
rect 35962 148934 36014 148986
rect 36066 148934 36118 148986
rect 66578 148934 66630 148986
rect 66682 148934 66734 148986
rect 66786 148934 66838 148986
rect 97298 148934 97350 148986
rect 97402 148934 97454 148986
rect 97506 148934 97558 148986
rect 128018 148934 128070 148986
rect 128122 148934 128174 148986
rect 128226 148934 128278 148986
rect 158738 148934 158790 148986
rect 158842 148934 158894 148986
rect 158946 148934 158998 148986
rect 189458 148934 189510 148986
rect 189562 148934 189614 148986
rect 189666 148934 189718 148986
rect 4478 148150 4530 148202
rect 4582 148150 4634 148202
rect 4686 148150 4738 148202
rect 35198 148150 35250 148202
rect 35302 148150 35354 148202
rect 35406 148150 35458 148202
rect 65918 148150 65970 148202
rect 66022 148150 66074 148202
rect 66126 148150 66178 148202
rect 96638 148150 96690 148202
rect 96742 148150 96794 148202
rect 96846 148150 96898 148202
rect 127358 148150 127410 148202
rect 127462 148150 127514 148202
rect 127566 148150 127618 148202
rect 158078 148150 158130 148202
rect 158182 148150 158234 148202
rect 158286 148150 158338 148202
rect 188798 148150 188850 148202
rect 188902 148150 188954 148202
rect 189006 148150 189058 148202
rect 5138 147366 5190 147418
rect 5242 147366 5294 147418
rect 5346 147366 5398 147418
rect 35858 147366 35910 147418
rect 35962 147366 36014 147418
rect 36066 147366 36118 147418
rect 66578 147366 66630 147418
rect 66682 147366 66734 147418
rect 66786 147366 66838 147418
rect 97298 147366 97350 147418
rect 97402 147366 97454 147418
rect 97506 147366 97558 147418
rect 128018 147366 128070 147418
rect 128122 147366 128174 147418
rect 128226 147366 128278 147418
rect 158738 147366 158790 147418
rect 158842 147366 158894 147418
rect 158946 147366 158998 147418
rect 189458 147366 189510 147418
rect 189562 147366 189614 147418
rect 189666 147366 189718 147418
rect 1822 146974 1874 147026
rect 2830 146862 2882 146914
rect 4478 146582 4530 146634
rect 4582 146582 4634 146634
rect 4686 146582 4738 146634
rect 35198 146582 35250 146634
rect 35302 146582 35354 146634
rect 35406 146582 35458 146634
rect 65918 146582 65970 146634
rect 66022 146582 66074 146634
rect 66126 146582 66178 146634
rect 96638 146582 96690 146634
rect 96742 146582 96794 146634
rect 96846 146582 96898 146634
rect 127358 146582 127410 146634
rect 127462 146582 127514 146634
rect 127566 146582 127618 146634
rect 158078 146582 158130 146634
rect 158182 146582 158234 146634
rect 158286 146582 158338 146634
rect 188798 146582 188850 146634
rect 188902 146582 188954 146634
rect 189006 146582 189058 146634
rect 1822 146302 1874 146354
rect 204094 146302 204146 146354
rect 201070 146190 201122 146242
rect 201742 146190 201794 146242
rect 5138 145798 5190 145850
rect 5242 145798 5294 145850
rect 5346 145798 5398 145850
rect 35858 145798 35910 145850
rect 35962 145798 36014 145850
rect 36066 145798 36118 145850
rect 66578 145798 66630 145850
rect 66682 145798 66734 145850
rect 66786 145798 66838 145850
rect 97298 145798 97350 145850
rect 97402 145798 97454 145850
rect 97506 145798 97558 145850
rect 128018 145798 128070 145850
rect 128122 145798 128174 145850
rect 128226 145798 128278 145850
rect 158738 145798 158790 145850
rect 158842 145798 158894 145850
rect 158946 145798 158998 145850
rect 189458 145798 189510 145850
rect 189562 145798 189614 145850
rect 189666 145798 189718 145850
rect 4478 145014 4530 145066
rect 4582 145014 4634 145066
rect 4686 145014 4738 145066
rect 35198 145014 35250 145066
rect 35302 145014 35354 145066
rect 35406 145014 35458 145066
rect 65918 145014 65970 145066
rect 66022 145014 66074 145066
rect 66126 145014 66178 145066
rect 96638 145014 96690 145066
rect 96742 145014 96794 145066
rect 96846 145014 96898 145066
rect 127358 145014 127410 145066
rect 127462 145014 127514 145066
rect 127566 145014 127618 145066
rect 158078 145014 158130 145066
rect 158182 145014 158234 145066
rect 158286 145014 158338 145066
rect 188798 145014 188850 145066
rect 188902 145014 188954 145066
rect 189006 145014 189058 145066
rect 5138 144230 5190 144282
rect 5242 144230 5294 144282
rect 5346 144230 5398 144282
rect 189458 144230 189510 144282
rect 189562 144230 189614 144282
rect 189666 144230 189718 144282
rect 4478 143446 4530 143498
rect 4582 143446 4634 143498
rect 4686 143446 4738 143498
rect 188798 143446 188850 143498
rect 188902 143446 188954 143498
rect 189006 143446 189058 143498
rect 1710 142830 1762 142882
rect 5138 142662 5190 142714
rect 5242 142662 5294 142714
rect 5346 142662 5398 142714
rect 189458 142662 189510 142714
rect 189562 142662 189614 142714
rect 189666 142662 189718 142714
rect 4478 141878 4530 141930
rect 4582 141878 4634 141930
rect 4686 141878 4738 141930
rect 188798 141878 188850 141930
rect 188902 141878 188954 141930
rect 189006 141878 189058 141930
rect 5138 141094 5190 141146
rect 5242 141094 5294 141146
rect 5346 141094 5398 141146
rect 189458 141094 189510 141146
rect 189562 141094 189614 141146
rect 189666 141094 189718 141146
rect 4478 140310 4530 140362
rect 4582 140310 4634 140362
rect 4686 140310 4738 140362
rect 188798 140310 188850 140362
rect 188902 140310 188954 140362
rect 189006 140310 189058 140362
rect 5138 139526 5190 139578
rect 5242 139526 5294 139578
rect 5346 139526 5398 139578
rect 189458 139526 189510 139578
rect 189562 139526 189614 139578
rect 189666 139526 189718 139578
rect 1710 138910 1762 138962
rect 4478 138742 4530 138794
rect 4582 138742 4634 138794
rect 4686 138742 4738 138794
rect 188798 138742 188850 138794
rect 188902 138742 188954 138794
rect 189006 138742 189058 138794
rect 5138 137958 5190 138010
rect 5242 137958 5294 138010
rect 5346 137958 5398 138010
rect 189458 137958 189510 138010
rect 189562 137958 189614 138010
rect 189666 137958 189718 138010
rect 4478 137174 4530 137226
rect 4582 137174 4634 137226
rect 4686 137174 4738 137226
rect 188798 137174 188850 137226
rect 188902 137174 188954 137226
rect 189006 137174 189058 137226
rect 5138 136390 5190 136442
rect 5242 136390 5294 136442
rect 5346 136390 5398 136442
rect 189458 136390 189510 136442
rect 189562 136390 189614 136442
rect 189666 136390 189718 136442
rect 4478 135606 4530 135658
rect 4582 135606 4634 135658
rect 4686 135606 4738 135658
rect 188798 135606 188850 135658
rect 188902 135606 188954 135658
rect 189006 135606 189058 135658
rect 1710 135214 1762 135266
rect 2830 135102 2882 135154
rect 5138 134822 5190 134874
rect 5242 134822 5294 134874
rect 5346 134822 5398 134874
rect 189458 134822 189510 134874
rect 189562 134822 189614 134874
rect 189666 134822 189718 134874
rect 1822 134654 1874 134706
rect 4478 134038 4530 134090
rect 4582 134038 4634 134090
rect 4686 134038 4738 134090
rect 188798 134038 188850 134090
rect 188902 134038 188954 134090
rect 189006 134038 189058 134090
rect 5138 133254 5190 133306
rect 5242 133254 5294 133306
rect 5346 133254 5398 133306
rect 189458 133254 189510 133306
rect 189562 133254 189614 133306
rect 189666 133254 189718 133306
rect 4478 132470 4530 132522
rect 4582 132470 4634 132522
rect 4686 132470 4738 132522
rect 188798 132470 188850 132522
rect 188902 132470 188954 132522
rect 189006 132470 189058 132522
rect 1710 131854 1762 131906
rect 5138 131686 5190 131738
rect 5242 131686 5294 131738
rect 5346 131686 5398 131738
rect 189458 131686 189510 131738
rect 189562 131686 189614 131738
rect 189666 131686 189718 131738
rect 4478 130902 4530 130954
rect 4582 130902 4634 130954
rect 4686 130902 4738 130954
rect 188798 130902 188850 130954
rect 188902 130902 188954 130954
rect 189006 130902 189058 130954
rect 5138 130118 5190 130170
rect 5242 130118 5294 130170
rect 5346 130118 5398 130170
rect 189458 130118 189510 130170
rect 189562 130118 189614 130170
rect 189666 130118 189718 130170
rect 4478 129334 4530 129386
rect 4582 129334 4634 129386
rect 4686 129334 4738 129386
rect 188798 129334 188850 129386
rect 188902 129334 188954 129386
rect 189006 129334 189058 129386
rect 5138 128550 5190 128602
rect 5242 128550 5294 128602
rect 5346 128550 5398 128602
rect 189458 128550 189510 128602
rect 189562 128550 189614 128602
rect 189666 128550 189718 128602
rect 203758 128270 203810 128322
rect 1710 127934 1762 127986
rect 4478 127766 4530 127818
rect 4582 127766 4634 127818
rect 4686 127766 4738 127818
rect 188798 127766 188850 127818
rect 188902 127766 188954 127818
rect 189006 127766 189058 127818
rect 5138 126982 5190 127034
rect 5242 126982 5294 127034
rect 5346 126982 5398 127034
rect 189458 126982 189510 127034
rect 189562 126982 189614 127034
rect 189666 126982 189718 127034
rect 4478 126198 4530 126250
rect 4582 126198 4634 126250
rect 4686 126198 4738 126250
rect 188798 126198 188850 126250
rect 188902 126198 188954 126250
rect 189006 126198 189058 126250
rect 5138 125414 5190 125466
rect 5242 125414 5294 125466
rect 5346 125414 5398 125466
rect 189458 125414 189510 125466
rect 189562 125414 189614 125466
rect 189666 125414 189718 125466
rect 4478 124630 4530 124682
rect 4582 124630 4634 124682
rect 4686 124630 4738 124682
rect 188798 124630 188850 124682
rect 188902 124630 188954 124682
rect 189006 124630 189058 124682
rect 1822 124238 1874 124290
rect 2830 124126 2882 124178
rect 5138 123846 5190 123898
rect 5242 123846 5294 123898
rect 5346 123846 5398 123898
rect 189458 123846 189510 123898
rect 189562 123846 189614 123898
rect 189666 123846 189718 123898
rect 1822 123678 1874 123730
rect 4478 123062 4530 123114
rect 4582 123062 4634 123114
rect 4686 123062 4738 123114
rect 188798 123062 188850 123114
rect 188902 123062 188954 123114
rect 189006 123062 189058 123114
rect 5138 122278 5190 122330
rect 5242 122278 5294 122330
rect 5346 122278 5398 122330
rect 189458 122278 189510 122330
rect 189562 122278 189614 122330
rect 189666 122278 189718 122330
rect 4478 121494 4530 121546
rect 4582 121494 4634 121546
rect 4686 121494 4738 121546
rect 188798 121494 188850 121546
rect 188902 121494 188954 121546
rect 189006 121494 189058 121546
rect 5138 120710 5190 120762
rect 5242 120710 5294 120762
rect 5346 120710 5398 120762
rect 189458 120710 189510 120762
rect 189562 120710 189614 120762
rect 189666 120710 189718 120762
rect 1710 120430 1762 120482
rect 4478 119926 4530 119978
rect 4582 119926 4634 119978
rect 4686 119926 4738 119978
rect 188798 119926 188850 119978
rect 188902 119926 188954 119978
rect 189006 119926 189058 119978
rect 204094 119646 204146 119698
rect 202190 119534 202242 119586
rect 5138 119142 5190 119194
rect 5242 119142 5294 119194
rect 5346 119142 5398 119194
rect 189458 119142 189510 119194
rect 189562 119142 189614 119194
rect 189666 119142 189718 119194
rect 203758 118638 203810 118690
rect 4478 118358 4530 118410
rect 4582 118358 4634 118410
rect 4686 118358 4738 118410
rect 188798 118358 188850 118410
rect 188902 118358 188954 118410
rect 189006 118358 189058 118410
rect 5138 117574 5190 117626
rect 5242 117574 5294 117626
rect 5346 117574 5398 117626
rect 189458 117574 189510 117626
rect 189562 117574 189614 117626
rect 189666 117574 189718 117626
rect 4478 116790 4530 116842
rect 4582 116790 4634 116842
rect 4686 116790 4738 116842
rect 188798 116790 188850 116842
rect 188902 116790 188954 116842
rect 189006 116790 189058 116842
rect 1710 116510 1762 116562
rect 5138 116006 5190 116058
rect 5242 116006 5294 116058
rect 5346 116006 5398 116058
rect 189458 116006 189510 116058
rect 189562 116006 189614 116058
rect 189666 116006 189718 116058
rect 4478 115222 4530 115274
rect 4582 115222 4634 115274
rect 4686 115222 4738 115274
rect 188798 115222 188850 115274
rect 188902 115222 188954 115274
rect 189006 115222 189058 115274
rect 5138 114438 5190 114490
rect 5242 114438 5294 114490
rect 5346 114438 5398 114490
rect 189458 114438 189510 114490
rect 189562 114438 189614 114490
rect 189666 114438 189718 114490
rect 4478 113654 4530 113706
rect 4582 113654 4634 113706
rect 4686 113654 4738 113706
rect 188798 113654 188850 113706
rect 188902 113654 188954 113706
rect 189006 113654 189058 113706
rect 5138 112870 5190 112922
rect 5242 112870 5294 112922
rect 5346 112870 5398 112922
rect 189458 112870 189510 112922
rect 189562 112870 189614 112922
rect 189666 112870 189718 112922
rect 1710 112478 1762 112530
rect 2830 112366 2882 112418
rect 4478 112086 4530 112138
rect 4582 112086 4634 112138
rect 4686 112086 4738 112138
rect 188798 112086 188850 112138
rect 188902 112086 188954 112138
rect 189006 112086 189058 112138
rect 1822 111806 1874 111858
rect 5138 111302 5190 111354
rect 5242 111302 5294 111354
rect 5346 111302 5398 111354
rect 189458 111302 189510 111354
rect 189562 111302 189614 111354
rect 189666 111302 189718 111354
rect 4478 110518 4530 110570
rect 4582 110518 4634 110570
rect 4686 110518 4738 110570
rect 188798 110518 188850 110570
rect 188902 110518 188954 110570
rect 189006 110518 189058 110570
rect 5138 109734 5190 109786
rect 5242 109734 5294 109786
rect 5346 109734 5398 109786
rect 189458 109734 189510 109786
rect 189562 109734 189614 109786
rect 189666 109734 189718 109786
rect 4478 108950 4530 109002
rect 4582 108950 4634 109002
rect 4686 108950 4738 109002
rect 188798 108950 188850 109002
rect 188902 108950 188954 109002
rect 189006 108950 189058 109002
rect 1710 108446 1762 108498
rect 5138 108166 5190 108218
rect 5242 108166 5294 108218
rect 5346 108166 5398 108218
rect 189458 108166 189510 108218
rect 189562 108166 189614 108218
rect 189666 108166 189718 108218
rect 4478 107382 4530 107434
rect 4582 107382 4634 107434
rect 4686 107382 4738 107434
rect 188798 107382 188850 107434
rect 188902 107382 188954 107434
rect 189006 107382 189058 107434
rect 5138 106598 5190 106650
rect 5242 106598 5294 106650
rect 5346 106598 5398 106650
rect 189458 106598 189510 106650
rect 189562 106598 189614 106650
rect 189666 106598 189718 106650
rect 4478 105814 4530 105866
rect 4582 105814 4634 105866
rect 4686 105814 4738 105866
rect 188798 105814 188850 105866
rect 188902 105814 188954 105866
rect 189006 105814 189058 105866
rect 1710 105534 1762 105586
rect 5138 105030 5190 105082
rect 5242 105030 5294 105082
rect 5346 105030 5398 105082
rect 189458 105030 189510 105082
rect 189562 105030 189614 105082
rect 189666 105030 189718 105082
rect 4478 104246 4530 104298
rect 4582 104246 4634 104298
rect 4686 104246 4738 104298
rect 188798 104246 188850 104298
rect 188902 104246 188954 104298
rect 189006 104246 189058 104298
rect 5138 103462 5190 103514
rect 5242 103462 5294 103514
rect 5346 103462 5398 103514
rect 189458 103462 189510 103514
rect 189562 103462 189614 103514
rect 189666 103462 189718 103514
rect 4478 102678 4530 102730
rect 4582 102678 4634 102730
rect 4686 102678 4738 102730
rect 188798 102678 188850 102730
rect 188902 102678 188954 102730
rect 189006 102678 189058 102730
rect 204318 102062 204370 102114
rect 5138 101894 5190 101946
rect 5242 101894 5294 101946
rect 5346 101894 5398 101946
rect 189458 101894 189510 101946
rect 189562 101894 189614 101946
rect 189666 101894 189718 101946
rect 2046 101614 2098 101666
rect 1710 101502 1762 101554
rect 2494 101390 2546 101442
rect 4478 101110 4530 101162
rect 4582 101110 4634 101162
rect 4686 101110 4738 101162
rect 188798 101110 188850 101162
rect 188902 101110 188954 101162
rect 189006 101110 189058 101162
rect 5138 100326 5190 100378
rect 5242 100326 5294 100378
rect 5346 100326 5398 100378
rect 189458 100326 189510 100378
rect 189562 100326 189614 100378
rect 189666 100326 189718 100378
rect 4478 99542 4530 99594
rect 4582 99542 4634 99594
rect 4686 99542 4738 99594
rect 188798 99542 188850 99594
rect 188902 99542 188954 99594
rect 189006 99542 189058 99594
rect 5138 98758 5190 98810
rect 5242 98758 5294 98810
rect 5346 98758 5398 98810
rect 189458 98758 189510 98810
rect 189562 98758 189614 98810
rect 189666 98758 189718 98810
rect 4478 97974 4530 98026
rect 4582 97974 4634 98026
rect 4686 97974 4738 98026
rect 188798 97974 188850 98026
rect 188902 97974 188954 98026
rect 189006 97974 189058 98026
rect 1710 97358 1762 97410
rect 5138 97190 5190 97242
rect 5242 97190 5294 97242
rect 5346 97190 5398 97242
rect 189458 97190 189510 97242
rect 189562 97190 189614 97242
rect 189666 97190 189718 97242
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 188798 96406 188850 96458
rect 188902 96406 188954 96458
rect 189006 96406 189058 96458
rect 5138 95622 5190 95674
rect 5242 95622 5294 95674
rect 5346 95622 5398 95674
rect 189458 95622 189510 95674
rect 189562 95622 189614 95674
rect 189666 95622 189718 95674
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 188798 94838 188850 94890
rect 188902 94838 188954 94890
rect 189006 94838 189058 94890
rect 5138 94054 5190 94106
rect 5242 94054 5294 94106
rect 5346 94054 5398 94106
rect 189458 94054 189510 94106
rect 189562 94054 189614 94106
rect 189666 94054 189718 94106
rect 201182 93662 201234 93714
rect 203198 93550 203250 93602
rect 1710 93438 1762 93490
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 188798 93270 188850 93322
rect 188902 93270 188954 93322
rect 189006 93270 189058 93322
rect 203982 92990 204034 93042
rect 5138 92486 5190 92538
rect 5242 92486 5294 92538
rect 5346 92486 5398 92538
rect 189458 92486 189510 92538
rect 189562 92486 189614 92538
rect 189666 92486 189718 92538
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 188798 91702 188850 91754
rect 188902 91702 188954 91754
rect 189006 91702 189058 91754
rect 5138 90918 5190 90970
rect 5242 90918 5294 90970
rect 5346 90918 5398 90970
rect 189458 90918 189510 90970
rect 189562 90918 189614 90970
rect 189666 90918 189718 90970
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 188798 90134 188850 90186
rect 188902 90134 188954 90186
rect 189006 90134 189058 90186
rect 1710 89518 1762 89570
rect 2046 89518 2098 89570
rect 2494 89518 2546 89570
rect 5138 89350 5190 89402
rect 5242 89350 5294 89402
rect 5346 89350 5398 89402
rect 189458 89350 189510 89402
rect 189562 89350 189614 89402
rect 189666 89350 189718 89402
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 188798 88566 188850 88618
rect 188902 88566 188954 88618
rect 189006 88566 189058 88618
rect 5138 87782 5190 87834
rect 5242 87782 5294 87834
rect 5346 87782 5398 87834
rect 189458 87782 189510 87834
rect 189562 87782 189614 87834
rect 189666 87782 189718 87834
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 188798 86998 188850 87050
rect 188902 86998 188954 87050
rect 189006 86998 189058 87050
rect 5138 86214 5190 86266
rect 5242 86214 5294 86266
rect 5346 86214 5398 86266
rect 189458 86214 189510 86266
rect 189562 86214 189614 86266
rect 189666 86214 189718 86266
rect 1710 85934 1762 85986
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 188798 85430 188850 85482
rect 188902 85430 188954 85482
rect 189006 85430 189058 85482
rect 5138 84646 5190 84698
rect 5242 84646 5294 84698
rect 5346 84646 5398 84698
rect 189458 84646 189510 84698
rect 189562 84646 189614 84698
rect 189666 84646 189718 84698
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 188798 83862 188850 83914
rect 188902 83862 188954 83914
rect 189006 83862 189058 83914
rect 5138 83078 5190 83130
rect 5242 83078 5294 83130
rect 5346 83078 5398 83130
rect 189458 83078 189510 83130
rect 189562 83078 189614 83130
rect 189666 83078 189718 83130
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 188798 82294 188850 82346
rect 188902 82294 188954 82346
rect 189006 82294 189058 82346
rect 1710 82014 1762 82066
rect 5138 81510 5190 81562
rect 5242 81510 5294 81562
rect 5346 81510 5398 81562
rect 189458 81510 189510 81562
rect 189562 81510 189614 81562
rect 189666 81510 189718 81562
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 188798 80726 188850 80778
rect 188902 80726 188954 80778
rect 189006 80726 189058 80778
rect 5138 79942 5190 79994
rect 5242 79942 5294 79994
rect 5346 79942 5398 79994
rect 189458 79942 189510 79994
rect 189562 79942 189614 79994
rect 189666 79942 189718 79994
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 188798 79158 188850 79210
rect 188902 79158 188954 79210
rect 189006 79158 189058 79210
rect 1710 78542 1762 78594
rect 2046 78542 2098 78594
rect 2494 78542 2546 78594
rect 17614 78542 17666 78594
rect 5138 78374 5190 78426
rect 5242 78374 5294 78426
rect 5346 78374 5398 78426
rect 189458 78374 189510 78426
rect 189562 78374 189614 78426
rect 189666 78374 189718 78426
rect 17614 77870 17666 77922
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 188798 77590 188850 77642
rect 188902 77590 188954 77642
rect 189006 77590 189058 77642
rect 5138 76806 5190 76858
rect 5242 76806 5294 76858
rect 5346 76806 5398 76858
rect 189458 76806 189510 76858
rect 189562 76806 189614 76858
rect 189666 76806 189718 76858
rect 17614 76302 17666 76354
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 188798 76022 188850 76074
rect 188902 76022 188954 76074
rect 189006 76022 189058 76074
rect 17502 75630 17554 75682
rect 204318 75518 204370 75570
rect 5138 75238 5190 75290
rect 5242 75238 5294 75290
rect 5346 75238 5398 75290
rect 189458 75238 189510 75290
rect 189562 75238 189614 75290
rect 189666 75238 189718 75290
rect 1710 74958 1762 75010
rect 17502 74734 17554 74786
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 188798 74454 188850 74506
rect 188902 74454 188954 74506
rect 189006 74454 189058 74506
rect 5138 73670 5190 73722
rect 5242 73670 5294 73722
rect 5346 73670 5398 73722
rect 189458 73670 189510 73722
rect 189562 73670 189614 73722
rect 189666 73670 189718 73722
rect 17502 73166 17554 73218
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 188798 72886 188850 72938
rect 188902 72886 188954 72938
rect 189006 72886 189058 72938
rect 5138 72102 5190 72154
rect 5242 72102 5294 72154
rect 5346 72102 5398 72154
rect 189458 72102 189510 72154
rect 189562 72102 189614 72154
rect 189666 72102 189718 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 188798 71318 188850 71370
rect 188902 71318 188954 71370
rect 189006 71318 189058 71370
rect 1710 71038 1762 71090
rect 5138 70534 5190 70586
rect 5242 70534 5294 70586
rect 5346 70534 5398 70586
rect 189458 70534 189510 70586
rect 189562 70534 189614 70586
rect 189666 70534 189718 70586
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 188798 69750 188850 69802
rect 188902 69750 188954 69802
rect 189006 69750 189058 69802
rect 5138 68966 5190 69018
rect 5242 68966 5294 69018
rect 5346 68966 5398 69018
rect 189458 68966 189510 69018
rect 189562 68966 189614 69018
rect 189666 68966 189718 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 188798 68182 188850 68234
rect 188902 68182 188954 68234
rect 189006 68182 189058 68234
rect 5138 67398 5190 67450
rect 5242 67398 5294 67450
rect 5346 67398 5398 67450
rect 189458 67398 189510 67450
rect 189562 67398 189614 67450
rect 189666 67398 189718 67450
rect 2046 67118 2098 67170
rect 1710 67006 1762 67058
rect 201182 67006 201234 67058
rect 2494 66894 2546 66946
rect 203198 66894 203250 66946
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 188798 66614 188850 66666
rect 188902 66614 188954 66666
rect 189006 66614 189058 66666
rect 203982 66334 204034 66386
rect 5138 65830 5190 65882
rect 5242 65830 5294 65882
rect 5346 65830 5398 65882
rect 189458 65830 189510 65882
rect 189562 65830 189614 65882
rect 189666 65830 189718 65882
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 188798 65046 188850 65098
rect 188902 65046 188954 65098
rect 189006 65046 189058 65098
rect 5138 64262 5190 64314
rect 5242 64262 5294 64314
rect 5346 64262 5398 64314
rect 189458 64262 189510 64314
rect 189562 64262 189614 64314
rect 189666 64262 189718 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 188798 63478 188850 63530
rect 188902 63478 188954 63530
rect 189006 63478 189058 63530
rect 1710 62862 1762 62914
rect 5138 62694 5190 62746
rect 5242 62694 5294 62746
rect 5346 62694 5398 62746
rect 189458 62694 189510 62746
rect 189562 62694 189614 62746
rect 189666 62694 189718 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 188798 61910 188850 61962
rect 188902 61910 188954 61962
rect 189006 61910 189058 61962
rect 5138 61126 5190 61178
rect 5242 61126 5294 61178
rect 5346 61126 5398 61178
rect 189458 61126 189510 61178
rect 189562 61126 189614 61178
rect 189666 61126 189718 61178
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 188798 60342 188850 60394
rect 188902 60342 188954 60394
rect 189006 60342 189058 60394
rect 5138 59558 5190 59610
rect 5242 59558 5294 59610
rect 5346 59558 5398 59610
rect 189458 59558 189510 59610
rect 189562 59558 189614 59610
rect 189666 59558 189718 59610
rect 1710 58942 1762 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 188798 58774 188850 58826
rect 188902 58774 188954 58826
rect 189006 58774 189058 58826
rect 5138 57990 5190 58042
rect 5242 57990 5294 58042
rect 5346 57990 5398 58042
rect 189458 57990 189510 58042
rect 189562 57990 189614 58042
rect 189666 57990 189718 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 188798 57206 188850 57258
rect 188902 57206 188954 57258
rect 189006 57206 189058 57258
rect 5138 56422 5190 56474
rect 5242 56422 5294 56474
rect 5346 56422 5398 56474
rect 189458 56422 189510 56474
rect 189562 56422 189614 56474
rect 189666 56422 189718 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 188798 55638 188850 55690
rect 188902 55638 188954 55690
rect 189006 55638 189058 55690
rect 2270 55246 2322 55298
rect 1710 55134 1762 55186
rect 5138 54854 5190 54906
rect 5242 54854 5294 54906
rect 5346 54854 5398 54906
rect 189458 54854 189510 54906
rect 189562 54854 189614 54906
rect 189666 54854 189718 54906
rect 1822 54686 1874 54738
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 188798 54070 188850 54122
rect 188902 54070 188954 54122
rect 189006 54070 189058 54122
rect 5138 53286 5190 53338
rect 5242 53286 5294 53338
rect 5346 53286 5398 53338
rect 189458 53286 189510 53338
rect 189562 53286 189614 53338
rect 189666 53286 189718 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 188798 52502 188850 52554
rect 188902 52502 188954 52554
rect 189006 52502 189058 52554
rect 1710 51886 1762 51938
rect 5138 51718 5190 51770
rect 5242 51718 5294 51770
rect 5346 51718 5398 51770
rect 189458 51718 189510 51770
rect 189562 51718 189614 51770
rect 189666 51718 189718 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 188798 50934 188850 50986
rect 188902 50934 188954 50986
rect 189006 50934 189058 50986
rect 5138 50150 5190 50202
rect 5242 50150 5294 50202
rect 5346 50150 5398 50202
rect 189458 50150 189510 50202
rect 189562 50150 189614 50202
rect 189666 50150 189718 50202
rect 203758 49870 203810 49922
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 188798 49366 188850 49418
rect 188902 49366 188954 49418
rect 189006 49366 189058 49418
rect 5138 48582 5190 48634
rect 5242 48582 5294 48634
rect 5346 48582 5398 48634
rect 189458 48582 189510 48634
rect 189562 48582 189614 48634
rect 189666 48582 189718 48634
rect 1710 47966 1762 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 188798 47798 188850 47850
rect 188902 47798 188954 47850
rect 189006 47798 189058 47850
rect 173966 47182 174018 47234
rect 174414 47182 174466 47234
rect 5138 47014 5190 47066
rect 5242 47014 5294 47066
rect 5346 47014 5398 47066
rect 189458 47014 189510 47066
rect 189562 47014 189614 47066
rect 189666 47014 189718 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 188798 46230 188850 46282
rect 188902 46230 188954 46282
rect 189006 46230 189058 46282
rect 5138 45446 5190 45498
rect 5242 45446 5294 45498
rect 5346 45446 5398 45498
rect 189458 45446 189510 45498
rect 189562 45446 189614 45498
rect 189666 45446 189718 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 188798 44662 188850 44714
rect 188902 44662 188954 44714
rect 189006 44662 189058 44714
rect 1822 44270 1874 44322
rect 2270 44270 2322 44322
rect 5138 43878 5190 43930
rect 5242 43878 5294 43930
rect 5346 43878 5398 43930
rect 189458 43878 189510 43930
rect 189562 43878 189614 43930
rect 189666 43878 189718 43930
rect 1822 43710 1874 43762
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 188798 43094 188850 43146
rect 188902 43094 188954 43146
rect 189006 43094 189058 43146
rect 5138 42310 5190 42362
rect 5242 42310 5294 42362
rect 5346 42310 5398 42362
rect 189458 42310 189510 42362
rect 189562 42310 189614 42362
rect 189666 42310 189718 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 188798 41526 188850 41578
rect 188902 41526 188954 41578
rect 189006 41526 189058 41578
rect 204094 41246 204146 41298
rect 201742 41134 201794 41186
rect 201406 40910 201458 40962
rect 5138 40742 5190 40794
rect 5242 40742 5294 40794
rect 5346 40742 5398 40794
rect 189458 40742 189510 40794
rect 189562 40742 189614 40794
rect 189666 40742 189718 40794
rect 1710 40462 1762 40514
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 188798 39958 188850 40010
rect 188902 39958 188954 40010
rect 189006 39958 189058 40010
rect 5138 39174 5190 39226
rect 5242 39174 5294 39226
rect 5346 39174 5398 39226
rect 189458 39174 189510 39226
rect 189562 39174 189614 39226
rect 189666 39174 189718 39226
rect 188750 38670 188802 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 188798 38390 188850 38442
rect 188902 38390 188954 38442
rect 189006 38390 189058 38442
rect 5138 37606 5190 37658
rect 5242 37606 5294 37658
rect 5346 37606 5398 37658
rect 189458 37606 189510 37658
rect 189562 37606 189614 37658
rect 189666 37606 189718 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 188798 36822 188850 36874
rect 188902 36822 188954 36874
rect 189006 36822 189058 36874
rect 1710 36542 1762 36594
rect 17614 36206 17666 36258
rect 5138 36038 5190 36090
rect 5242 36038 5294 36090
rect 5346 36038 5398 36090
rect 189458 36038 189510 36090
rect 189562 36038 189614 36090
rect 189666 36038 189718 36090
rect 16942 35534 16994 35586
rect 17614 35534 17666 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 188798 35254 188850 35306
rect 188902 35254 188954 35306
rect 189006 35254 189058 35306
rect 5138 34470 5190 34522
rect 5242 34470 5294 34522
rect 5346 34470 5398 34522
rect 189458 34470 189510 34522
rect 189562 34470 189614 34522
rect 189666 34470 189718 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 188798 33686 188850 33738
rect 188902 33686 188954 33738
rect 189006 33686 189058 33738
rect 5138 32902 5190 32954
rect 5242 32902 5294 32954
rect 5346 32902 5398 32954
rect 189458 32902 189510 32954
rect 189562 32902 189614 32954
rect 189666 32902 189718 32954
rect 2046 32734 2098 32786
rect 1710 32510 1762 32562
rect 2494 32398 2546 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 188798 32118 188850 32170
rect 188902 32118 188954 32170
rect 189006 32118 189058 32170
rect 5138 31334 5190 31386
rect 5242 31334 5294 31386
rect 5346 31334 5398 31386
rect 189458 31334 189510 31386
rect 189562 31334 189614 31386
rect 189666 31334 189718 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 188798 30550 188850 30602
rect 188902 30550 188954 30602
rect 189006 30550 189058 30602
rect 5138 29766 5190 29818
rect 5242 29766 5294 29818
rect 5346 29766 5398 29818
rect 189458 29766 189510 29818
rect 189562 29766 189614 29818
rect 189666 29766 189718 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 188798 28982 188850 29034
rect 188902 28982 188954 29034
rect 189006 28982 189058 29034
rect 1710 28478 1762 28530
rect 5138 28198 5190 28250
rect 5242 28198 5294 28250
rect 5346 28198 5398 28250
rect 189458 28198 189510 28250
rect 189562 28198 189614 28250
rect 189666 28198 189718 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 188798 27414 188850 27466
rect 188902 27414 188954 27466
rect 189006 27414 189058 27466
rect 5138 26630 5190 26682
rect 5242 26630 5294 26682
rect 5346 26630 5398 26682
rect 189458 26630 189510 26682
rect 189562 26630 189614 26682
rect 189666 26630 189718 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 188798 25846 188850 25898
rect 188902 25846 188954 25898
rect 189006 25846 189058 25898
rect 1710 25566 1762 25618
rect 5138 25062 5190 25114
rect 5242 25062 5294 25114
rect 5346 25062 5398 25114
rect 189458 25062 189510 25114
rect 189562 25062 189614 25114
rect 189666 25062 189718 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 188798 24278 188850 24330
rect 188902 24278 188954 24330
rect 189006 24278 189058 24330
rect 204318 23662 204370 23714
rect 5138 23494 5190 23546
rect 5242 23494 5294 23546
rect 5346 23494 5398 23546
rect 189458 23494 189510 23546
rect 189562 23494 189614 23546
rect 189666 23494 189718 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 188798 22710 188850 22762
rect 188902 22710 188954 22762
rect 189006 22710 189058 22762
rect 5138 21926 5190 21978
rect 5242 21926 5294 21978
rect 5346 21926 5398 21978
rect 189458 21926 189510 21978
rect 189562 21926 189614 21978
rect 189666 21926 189718 21978
rect 2046 21758 2098 21810
rect 1710 21534 1762 21586
rect 2494 21422 2546 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 188798 21142 188850 21194
rect 188902 21142 188954 21194
rect 189006 21142 189058 21194
rect 5138 20358 5190 20410
rect 5242 20358 5294 20410
rect 5346 20358 5398 20410
rect 189458 20358 189510 20410
rect 189562 20358 189614 20410
rect 189666 20358 189718 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 188798 19574 188850 19626
rect 188902 19574 188954 19626
rect 189006 19574 189058 19626
rect 5138 18790 5190 18842
rect 5242 18790 5294 18842
rect 5346 18790 5398 18842
rect 189458 18790 189510 18842
rect 189562 18790 189614 18842
rect 189666 18790 189718 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 188798 18006 188850 18058
rect 188902 18006 188954 18058
rect 189006 18006 189058 18058
rect 1710 17390 1762 17442
rect 5138 17222 5190 17274
rect 5242 17222 5294 17274
rect 5346 17222 5398 17274
rect 35858 17222 35910 17274
rect 35962 17222 36014 17274
rect 36066 17222 36118 17274
rect 66578 17222 66630 17274
rect 66682 17222 66734 17274
rect 66786 17222 66838 17274
rect 97298 17222 97350 17274
rect 97402 17222 97454 17274
rect 97506 17222 97558 17274
rect 128018 17222 128070 17274
rect 128122 17222 128174 17274
rect 128226 17222 128278 17274
rect 158738 17222 158790 17274
rect 158842 17222 158894 17274
rect 158946 17222 158998 17274
rect 189458 17222 189510 17274
rect 189562 17222 189614 17274
rect 189666 17222 189718 17274
rect 44718 17054 44770 17106
rect 48190 17054 48242 17106
rect 51550 17054 51602 17106
rect 55134 17054 55186 17106
rect 59054 17054 59106 17106
rect 61966 17054 62018 17106
rect 65438 17054 65490 17106
rect 68798 17054 68850 17106
rect 72158 17054 72210 17106
rect 75518 17054 75570 17106
rect 78990 17054 79042 17106
rect 82350 17054 82402 17106
rect 82910 17054 82962 17106
rect 97134 17054 97186 17106
rect 111246 17054 111298 17106
rect 140030 17054 140082 17106
rect 154366 17054 154418 17106
rect 67902 16830 67954 16882
rect 125582 16830 125634 16882
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 127358 16438 127410 16490
rect 127462 16438 127514 16490
rect 127566 16438 127618 16490
rect 158078 16438 158130 16490
rect 158182 16438 158234 16490
rect 158286 16438 158338 16490
rect 188798 16438 188850 16490
rect 188902 16438 188954 16490
rect 189006 16438 189058 16490
rect 5138 15654 5190 15706
rect 5242 15654 5294 15706
rect 5346 15654 5398 15706
rect 35858 15654 35910 15706
rect 35962 15654 36014 15706
rect 36066 15654 36118 15706
rect 66578 15654 66630 15706
rect 66682 15654 66734 15706
rect 66786 15654 66838 15706
rect 97298 15654 97350 15706
rect 97402 15654 97454 15706
rect 97506 15654 97558 15706
rect 128018 15654 128070 15706
rect 128122 15654 128174 15706
rect 128226 15654 128278 15706
rect 158738 15654 158790 15706
rect 158842 15654 158894 15706
rect 158946 15654 158998 15706
rect 189458 15654 189510 15706
rect 189562 15654 189614 15706
rect 189666 15654 189718 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 127358 14870 127410 14922
rect 127462 14870 127514 14922
rect 127566 14870 127618 14922
rect 158078 14870 158130 14922
rect 158182 14870 158234 14922
rect 158286 14870 158338 14922
rect 188798 14870 188850 14922
rect 188902 14870 188954 14922
rect 189006 14870 189058 14922
rect 204094 14590 204146 14642
rect 201742 14478 201794 14530
rect 5138 14086 5190 14138
rect 5242 14086 5294 14138
rect 5346 14086 5398 14138
rect 35858 14086 35910 14138
rect 35962 14086 36014 14138
rect 36066 14086 36118 14138
rect 66578 14086 66630 14138
rect 66682 14086 66734 14138
rect 66786 14086 66838 14138
rect 97298 14086 97350 14138
rect 97402 14086 97454 14138
rect 97506 14086 97558 14138
rect 128018 14086 128070 14138
rect 128122 14086 128174 14138
rect 128226 14086 128278 14138
rect 158738 14086 158790 14138
rect 158842 14086 158894 14138
rect 158946 14086 158998 14138
rect 189458 14086 189510 14138
rect 189562 14086 189614 14138
rect 189666 14086 189718 14138
rect 204318 13918 204370 13970
rect 1710 13470 1762 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 127358 13302 127410 13354
rect 127462 13302 127514 13354
rect 127566 13302 127618 13354
rect 158078 13302 158130 13354
rect 158182 13302 158234 13354
rect 158286 13302 158338 13354
rect 188798 13302 188850 13354
rect 188902 13302 188954 13354
rect 189006 13302 189058 13354
rect 5138 12518 5190 12570
rect 5242 12518 5294 12570
rect 5346 12518 5398 12570
rect 35858 12518 35910 12570
rect 35962 12518 36014 12570
rect 36066 12518 36118 12570
rect 66578 12518 66630 12570
rect 66682 12518 66734 12570
rect 66786 12518 66838 12570
rect 97298 12518 97350 12570
rect 97402 12518 97454 12570
rect 97506 12518 97558 12570
rect 128018 12518 128070 12570
rect 128122 12518 128174 12570
rect 128226 12518 128278 12570
rect 158738 12518 158790 12570
rect 158842 12518 158894 12570
rect 158946 12518 158998 12570
rect 189458 12518 189510 12570
rect 189562 12518 189614 12570
rect 189666 12518 189718 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 127358 11734 127410 11786
rect 127462 11734 127514 11786
rect 127566 11734 127618 11786
rect 158078 11734 158130 11786
rect 158182 11734 158234 11786
rect 158286 11734 158338 11786
rect 188798 11734 188850 11786
rect 188902 11734 188954 11786
rect 189006 11734 189058 11786
rect 5138 10950 5190 11002
rect 5242 10950 5294 11002
rect 5346 10950 5398 11002
rect 35858 10950 35910 11002
rect 35962 10950 36014 11002
rect 36066 10950 36118 11002
rect 66578 10950 66630 11002
rect 66682 10950 66734 11002
rect 66786 10950 66838 11002
rect 97298 10950 97350 11002
rect 97402 10950 97454 11002
rect 97506 10950 97558 11002
rect 128018 10950 128070 11002
rect 128122 10950 128174 11002
rect 128226 10950 128278 11002
rect 158738 10950 158790 11002
rect 158842 10950 158894 11002
rect 158946 10950 158998 11002
rect 189458 10950 189510 11002
rect 189562 10950 189614 11002
rect 189666 10950 189718 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 127358 10166 127410 10218
rect 127462 10166 127514 10218
rect 127566 10166 127618 10218
rect 158078 10166 158130 10218
rect 158182 10166 158234 10218
rect 158286 10166 158338 10218
rect 188798 10166 188850 10218
rect 188902 10166 188954 10218
rect 189006 10166 189058 10218
rect 1710 9550 1762 9602
rect 2046 9550 2098 9602
rect 2494 9550 2546 9602
rect 5138 9382 5190 9434
rect 5242 9382 5294 9434
rect 5346 9382 5398 9434
rect 35858 9382 35910 9434
rect 35962 9382 36014 9434
rect 36066 9382 36118 9434
rect 66578 9382 66630 9434
rect 66682 9382 66734 9434
rect 66786 9382 66838 9434
rect 97298 9382 97350 9434
rect 97402 9382 97454 9434
rect 97506 9382 97558 9434
rect 128018 9382 128070 9434
rect 128122 9382 128174 9434
rect 128226 9382 128278 9434
rect 158738 9382 158790 9434
rect 158842 9382 158894 9434
rect 158946 9382 158998 9434
rect 189458 9382 189510 9434
rect 189562 9382 189614 9434
rect 189666 9382 189718 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 127358 8598 127410 8650
rect 127462 8598 127514 8650
rect 127566 8598 127618 8650
rect 158078 8598 158130 8650
rect 158182 8598 158234 8650
rect 158286 8598 158338 8650
rect 188798 8598 188850 8650
rect 188902 8598 188954 8650
rect 189006 8598 189058 8650
rect 5138 7814 5190 7866
rect 5242 7814 5294 7866
rect 5346 7814 5398 7866
rect 35858 7814 35910 7866
rect 35962 7814 36014 7866
rect 36066 7814 36118 7866
rect 66578 7814 66630 7866
rect 66682 7814 66734 7866
rect 66786 7814 66838 7866
rect 97298 7814 97350 7866
rect 97402 7814 97454 7866
rect 97506 7814 97558 7866
rect 128018 7814 128070 7866
rect 128122 7814 128174 7866
rect 128226 7814 128278 7866
rect 158738 7814 158790 7866
rect 158842 7814 158894 7866
rect 158946 7814 158998 7866
rect 189458 7814 189510 7866
rect 189562 7814 189614 7866
rect 189666 7814 189718 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 127358 7030 127410 7082
rect 127462 7030 127514 7082
rect 127566 7030 127618 7082
rect 158078 7030 158130 7082
rect 158182 7030 158234 7082
rect 158286 7030 158338 7082
rect 188798 7030 188850 7082
rect 188902 7030 188954 7082
rect 189006 7030 189058 7082
rect 5138 6246 5190 6298
rect 5242 6246 5294 6298
rect 5346 6246 5398 6298
rect 35858 6246 35910 6298
rect 35962 6246 36014 6298
rect 36066 6246 36118 6298
rect 66578 6246 66630 6298
rect 66682 6246 66734 6298
rect 66786 6246 66838 6298
rect 97298 6246 97350 6298
rect 97402 6246 97454 6298
rect 97506 6246 97558 6298
rect 128018 6246 128070 6298
rect 128122 6246 128174 6298
rect 128226 6246 128278 6298
rect 158738 6246 158790 6298
rect 158842 6246 158894 6298
rect 158946 6246 158998 6298
rect 189458 6246 189510 6298
rect 189562 6246 189614 6298
rect 189666 6246 189718 6298
rect 1710 5966 1762 6018
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 127358 5462 127410 5514
rect 127462 5462 127514 5514
rect 127566 5462 127618 5514
rect 158078 5462 158130 5514
rect 158182 5462 158234 5514
rect 158286 5462 158338 5514
rect 188798 5462 188850 5514
rect 188902 5462 188954 5514
rect 189006 5462 189058 5514
rect 5138 4678 5190 4730
rect 5242 4678 5294 4730
rect 5346 4678 5398 4730
rect 35858 4678 35910 4730
rect 35962 4678 36014 4730
rect 36066 4678 36118 4730
rect 66578 4678 66630 4730
rect 66682 4678 66734 4730
rect 66786 4678 66838 4730
rect 97298 4678 97350 4730
rect 97402 4678 97454 4730
rect 97506 4678 97558 4730
rect 128018 4678 128070 4730
rect 128122 4678 128174 4730
rect 128226 4678 128278 4730
rect 158738 4678 158790 4730
rect 158842 4678 158894 4730
rect 158946 4678 158998 4730
rect 189458 4678 189510 4730
rect 189562 4678 189614 4730
rect 189666 4678 189718 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 127358 3894 127410 3946
rect 127462 3894 127514 3946
rect 127566 3894 127618 3946
rect 158078 3894 158130 3946
rect 158182 3894 158234 3946
rect 158286 3894 158338 3946
rect 188798 3894 188850 3946
rect 188902 3894 188954 3946
rect 189006 3894 189058 3946
rect 1710 3614 1762 3666
rect 34526 3278 34578 3330
rect 103070 3278 103122 3330
rect 171614 3278 171666 3330
rect 5138 3110 5190 3162
rect 5242 3110 5294 3162
rect 5346 3110 5398 3162
rect 35858 3110 35910 3162
rect 35962 3110 36014 3162
rect 36066 3110 36118 3162
rect 66578 3110 66630 3162
rect 66682 3110 66734 3162
rect 66786 3110 66838 3162
rect 97298 3110 97350 3162
rect 97402 3110 97454 3162
rect 97506 3110 97558 3162
rect 128018 3110 128070 3162
rect 128122 3110 128174 3162
rect 128226 3110 128278 3162
rect 158738 3110 158790 3162
rect 158842 3110 158894 3162
rect 158946 3110 158998 3162
rect 189458 3110 189510 3162
rect 189562 3110 189614 3162
rect 189666 3110 189718 3162
<< metal2 >>
rect 3808 159264 3920 160064
rect 11424 159264 11536 160064
rect 19040 159264 19152 160064
rect 26656 159264 26768 160064
rect 34272 159264 34384 160064
rect 41888 159264 42000 160064
rect 49504 159264 49616 160064
rect 57120 159264 57232 160064
rect 64736 159264 64848 160064
rect 72352 159264 72464 160064
rect 79968 159264 80080 160064
rect 87584 159264 87696 160064
rect 95200 159264 95312 160064
rect 102816 159264 102928 160064
rect 110432 159264 110544 160064
rect 118048 159264 118160 160064
rect 125664 159264 125776 160064
rect 133280 159264 133392 160064
rect 140896 159264 141008 160064
rect 148512 159264 148624 160064
rect 156128 159264 156240 160064
rect 163744 159264 163856 160064
rect 171360 159264 171472 160064
rect 178976 159264 179088 160064
rect 186592 159264 186704 160064
rect 194208 159264 194320 160064
rect 201824 159264 201936 160064
rect 1708 157892 1764 157902
rect 1708 156548 1764 157836
rect 1708 156546 1876 156548
rect 1708 156494 1710 156546
rect 1762 156494 1876 156546
rect 1708 156492 1876 156494
rect 1708 156482 1764 156492
rect 1820 155762 1876 156492
rect 1820 155710 1822 155762
rect 1874 155710 1876 155762
rect 1820 155698 1876 155710
rect 2380 156322 2436 156334
rect 2380 156270 2382 156322
rect 2434 156270 2436 156322
rect 1708 154978 1764 154990
rect 1708 154926 1710 154978
rect 1762 154926 1764 154978
rect 1708 154196 1764 154926
rect 1708 154130 1764 154140
rect 1708 151058 1764 151070
rect 1708 151006 1710 151058
rect 1762 151006 1764 151058
rect 1708 150388 1764 151006
rect 1708 150322 1764 150332
rect 1820 147026 1876 147038
rect 1820 146974 1822 147026
rect 1874 146974 1876 147026
rect 1820 146580 1876 146974
rect 1820 146354 1876 146524
rect 1820 146302 1822 146354
rect 1874 146302 1876 146354
rect 1820 146290 1876 146302
rect 1708 142882 1764 142894
rect 1708 142830 1710 142882
rect 1762 142830 1764 142882
rect 1708 142772 1764 142830
rect 1708 142706 1764 142716
rect 1708 138964 1764 138974
rect 1708 138870 1764 138908
rect 1708 135266 1764 135278
rect 1708 135214 1710 135266
rect 1762 135214 1764 135266
rect 1708 135156 1764 135214
rect 1708 134708 1764 135100
rect 1820 134708 1876 134718
rect 1708 134706 1876 134708
rect 1708 134654 1822 134706
rect 1874 134654 1876 134706
rect 1708 134652 1876 134654
rect 1820 134642 1876 134652
rect 1708 131906 1764 131918
rect 1708 131854 1710 131906
rect 1762 131854 1764 131906
rect 1708 131348 1764 131854
rect 1708 131282 1764 131292
rect 1708 127986 1764 127998
rect 1708 127934 1710 127986
rect 1762 127934 1764 127986
rect 1708 127540 1764 127934
rect 1708 127474 1764 127484
rect 1820 124290 1876 124302
rect 1820 124238 1822 124290
rect 1874 124238 1876 124290
rect 1820 123732 1876 124238
rect 1820 123638 1876 123676
rect 1708 120482 1764 120494
rect 1708 120430 1710 120482
rect 1762 120430 1764 120482
rect 1708 119924 1764 120430
rect 1708 119858 1764 119868
rect 1708 116562 1764 116574
rect 1708 116510 1710 116562
rect 1762 116510 1764 116562
rect 1708 116116 1764 116510
rect 1708 116050 1764 116060
rect 1708 112530 1764 112542
rect 1708 112478 1710 112530
rect 1762 112478 1764 112530
rect 1708 112308 1764 112478
rect 1764 112252 1876 112308
rect 1708 112242 1764 112252
rect 1820 111858 1876 112252
rect 1820 111806 1822 111858
rect 1874 111806 1876 111858
rect 1820 111794 1876 111806
rect 1708 108500 1764 108510
rect 1708 108406 1764 108444
rect 1708 105586 1764 105598
rect 1708 105534 1710 105586
rect 1762 105534 1764 105586
rect 1708 104692 1764 105534
rect 1708 104626 1764 104636
rect 2044 101668 2100 101678
rect 2044 101574 2100 101612
rect 1708 101554 1764 101566
rect 1708 101502 1710 101554
rect 1762 101502 1764 101554
rect 1708 101444 1764 101502
rect 1708 100884 1764 101388
rect 1708 100818 1764 100828
rect 1708 97410 1764 97422
rect 1708 97358 1710 97410
rect 1762 97358 1764 97410
rect 1708 97076 1764 97358
rect 1708 97010 1764 97020
rect 1708 93492 1764 93502
rect 1708 93398 1764 93436
rect 1708 89570 1764 89582
rect 1708 89518 1710 89570
rect 1762 89518 1764 89570
rect 1708 89460 1764 89518
rect 1708 89394 1764 89404
rect 2044 89570 2100 89582
rect 2044 89518 2046 89570
rect 2098 89518 2100 89570
rect 1708 85986 1764 85998
rect 1708 85934 1710 85986
rect 1762 85934 1764 85986
rect 1708 85652 1764 85934
rect 1708 85586 1764 85596
rect 1708 82068 1764 82078
rect 1708 81974 1764 82012
rect 2044 78988 2100 89518
rect 2044 78932 2212 78988
rect 1708 78596 1764 78606
rect 1708 78036 1764 78540
rect 1708 77970 1764 77980
rect 2044 78594 2100 78606
rect 2044 78542 2046 78594
rect 2098 78542 2100 78594
rect 2044 75684 2100 78542
rect 2044 75618 2100 75628
rect 1708 75010 1764 75022
rect 1708 74958 1710 75010
rect 1762 74958 1764 75010
rect 1708 74228 1764 74958
rect 2156 74788 2212 78932
rect 2156 74722 2212 74732
rect 2268 76356 2324 76366
rect 1708 74162 1764 74172
rect 1708 71090 1764 71102
rect 1708 71038 1710 71090
rect 1762 71038 1764 71090
rect 1708 70420 1764 71038
rect 1708 70354 1764 70364
rect 2268 67228 2324 76300
rect 2044 67172 2324 67228
rect 2044 67170 2100 67172
rect 2044 67118 2046 67170
rect 2098 67118 2100 67170
rect 2044 67106 2100 67118
rect 1708 67058 1764 67070
rect 1708 67006 1710 67058
rect 1762 67006 1764 67058
rect 1708 66612 1764 67006
rect 1708 66546 1764 66556
rect 1708 62916 1764 62926
rect 1708 62822 1764 62860
rect 1708 58996 1764 59006
rect 1708 58902 1764 58940
rect 2268 55300 2324 55310
rect 2268 55206 2324 55244
rect 1708 55188 1764 55198
rect 1708 54740 1764 55132
rect 1820 54740 1876 54750
rect 1708 54738 1876 54740
rect 1708 54686 1822 54738
rect 1874 54686 1876 54738
rect 1708 54684 1876 54686
rect 1820 54674 1876 54684
rect 1708 51938 1764 51950
rect 1708 51886 1710 51938
rect 1762 51886 1764 51938
rect 1708 51380 1764 51886
rect 1708 51314 1764 51324
rect 1708 48018 1764 48030
rect 1708 47966 1710 48018
rect 1762 47966 1764 48018
rect 1708 47572 1764 47966
rect 1708 47506 1764 47516
rect 1820 44322 1876 44334
rect 1820 44270 1822 44322
rect 1874 44270 1876 44322
rect 1820 43764 1876 44270
rect 2268 44324 2324 44334
rect 2268 44230 2324 44268
rect 1820 43698 1876 43708
rect 1708 40514 1764 40526
rect 1708 40462 1710 40514
rect 1762 40462 1764 40514
rect 1708 39956 1764 40462
rect 1708 39890 1764 39900
rect 1708 36594 1764 36606
rect 1708 36542 1710 36594
rect 1762 36542 1764 36594
rect 1708 36148 1764 36542
rect 1708 36082 1764 36092
rect 2044 36260 2100 36270
rect 2044 32786 2100 36204
rect 2044 32734 2046 32786
rect 2098 32734 2100 32786
rect 2044 32722 2100 32734
rect 2156 34692 2212 34702
rect 1708 32562 1764 32574
rect 1708 32510 1710 32562
rect 1762 32510 1764 32562
rect 1708 32340 1764 32510
rect 1708 32274 1764 32284
rect 1708 28532 1764 28542
rect 1708 28438 1764 28476
rect 1708 25618 1764 25630
rect 1708 25566 1710 25618
rect 1762 25566 1764 25618
rect 1708 24724 1764 25566
rect 1708 24658 1764 24668
rect 2044 21812 2100 21822
rect 2156 21812 2212 34636
rect 2380 29428 2436 156270
rect 3836 156212 3892 159264
rect 5136 156828 5400 156838
rect 5192 156772 5240 156828
rect 5296 156772 5344 156828
rect 5136 156762 5400 156772
rect 11452 156660 11508 159264
rect 11676 156660 11732 156670
rect 11452 156658 11732 156660
rect 11452 156606 11678 156658
rect 11730 156606 11732 156658
rect 11452 156604 11732 156606
rect 11676 156594 11732 156604
rect 19068 156660 19124 159264
rect 19292 156660 19348 156670
rect 19068 156658 19348 156660
rect 19068 156606 19070 156658
rect 19122 156606 19294 156658
rect 19346 156606 19348 156658
rect 19068 156604 19348 156606
rect 19068 156594 19124 156604
rect 19292 156594 19348 156604
rect 20076 156324 20132 156334
rect 20076 156230 20132 156268
rect 22764 156324 22820 156334
rect 4060 156212 4116 156222
rect 3836 156210 4116 156212
rect 3836 156158 4062 156210
rect 4114 156158 4116 156210
rect 3836 156156 4116 156158
rect 4060 156146 4116 156156
rect 4476 156044 4740 156054
rect 4532 155988 4580 156044
rect 4636 155988 4684 156044
rect 4476 155978 4740 155988
rect 5136 155260 5400 155270
rect 5192 155204 5240 155260
rect 5296 155204 5344 155260
rect 5136 155194 5400 155204
rect 4476 154476 4740 154486
rect 4532 154420 4580 154476
rect 4636 154420 4684 154476
rect 4476 154410 4740 154420
rect 5136 153692 5400 153702
rect 5192 153636 5240 153692
rect 5296 153636 5344 153692
rect 5136 153626 5400 153636
rect 4476 152908 4740 152918
rect 4532 152852 4580 152908
rect 4636 152852 4684 152908
rect 4476 152842 4740 152852
rect 5136 152124 5400 152134
rect 5192 152068 5240 152124
rect 5296 152068 5344 152124
rect 5136 152058 5400 152068
rect 4476 151340 4740 151350
rect 4532 151284 4580 151340
rect 4636 151284 4684 151340
rect 4476 151274 4740 151284
rect 5136 150556 5400 150566
rect 5192 150500 5240 150556
rect 5296 150500 5344 150556
rect 5136 150490 5400 150500
rect 4476 149772 4740 149782
rect 4532 149716 4580 149772
rect 4636 149716 4684 149772
rect 4476 149706 4740 149716
rect 5136 148988 5400 148998
rect 5192 148932 5240 148988
rect 5296 148932 5344 148988
rect 5136 148922 5400 148932
rect 4476 148204 4740 148214
rect 4532 148148 4580 148204
rect 4636 148148 4684 148204
rect 4476 148138 4740 148148
rect 5136 147420 5400 147430
rect 5192 147364 5240 147420
rect 5296 147364 5344 147420
rect 5136 147354 5400 147364
rect 2828 146916 2884 146926
rect 2828 146822 2884 146860
rect 12572 146916 12628 146926
rect 4476 146636 4740 146646
rect 4532 146580 4580 146636
rect 4636 146580 4684 146636
rect 4476 146570 4740 146580
rect 5136 145852 5400 145862
rect 5192 145796 5240 145852
rect 5296 145796 5344 145852
rect 5136 145786 5400 145796
rect 4476 145068 4740 145078
rect 4532 145012 4580 145068
rect 4636 145012 4684 145068
rect 4476 145002 4740 145012
rect 5136 144284 5400 144294
rect 5192 144228 5240 144284
rect 5296 144228 5344 144284
rect 5136 144218 5400 144228
rect 4476 143500 4740 143510
rect 4532 143444 4580 143500
rect 4636 143444 4684 143500
rect 4476 143434 4740 143444
rect 5136 142716 5400 142726
rect 5192 142660 5240 142716
rect 5296 142660 5344 142716
rect 5136 142650 5400 142660
rect 4476 141932 4740 141942
rect 4532 141876 4580 141932
rect 4636 141876 4684 141932
rect 4476 141866 4740 141876
rect 5136 141148 5400 141158
rect 5192 141092 5240 141148
rect 5296 141092 5344 141148
rect 5136 141082 5400 141092
rect 4476 140364 4740 140374
rect 4532 140308 4580 140364
rect 4636 140308 4684 140364
rect 4476 140298 4740 140308
rect 5136 139580 5400 139590
rect 5192 139524 5240 139580
rect 5296 139524 5344 139580
rect 5136 139514 5400 139524
rect 4476 138796 4740 138806
rect 4532 138740 4580 138796
rect 4636 138740 4684 138796
rect 4476 138730 4740 138740
rect 5136 138012 5400 138022
rect 5192 137956 5240 138012
rect 5296 137956 5344 138012
rect 5136 137946 5400 137956
rect 4476 137228 4740 137238
rect 4532 137172 4580 137228
rect 4636 137172 4684 137228
rect 4476 137162 4740 137172
rect 5136 136444 5400 136454
rect 5192 136388 5240 136444
rect 5296 136388 5344 136444
rect 5136 136378 5400 136388
rect 4476 135660 4740 135670
rect 4532 135604 4580 135660
rect 4636 135604 4684 135660
rect 4476 135594 4740 135604
rect 2828 135156 2884 135166
rect 2828 135062 2884 135100
rect 5136 134876 5400 134886
rect 5192 134820 5240 134876
rect 5296 134820 5344 134876
rect 5136 134810 5400 134820
rect 4476 134092 4740 134102
rect 4532 134036 4580 134092
rect 4636 134036 4684 134092
rect 4476 134026 4740 134036
rect 5136 133308 5400 133318
rect 5192 133252 5240 133308
rect 5296 133252 5344 133308
rect 5136 133242 5400 133252
rect 4476 132524 4740 132534
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4476 132458 4740 132468
rect 5136 131740 5400 131750
rect 5192 131684 5240 131740
rect 5296 131684 5344 131740
rect 5136 131674 5400 131684
rect 4476 130956 4740 130966
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4476 130890 4740 130900
rect 5136 130172 5400 130182
rect 5192 130116 5240 130172
rect 5296 130116 5344 130172
rect 5136 130106 5400 130116
rect 4476 129388 4740 129398
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4476 129322 4740 129332
rect 5136 128604 5400 128614
rect 5192 128548 5240 128604
rect 5296 128548 5344 128604
rect 5136 128538 5400 128548
rect 4476 127820 4740 127830
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4476 127754 4740 127764
rect 5136 127036 5400 127046
rect 5192 126980 5240 127036
rect 5296 126980 5344 127036
rect 5136 126970 5400 126980
rect 4476 126252 4740 126262
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4476 126186 4740 126196
rect 5136 125468 5400 125478
rect 5192 125412 5240 125468
rect 5296 125412 5344 125468
rect 5136 125402 5400 125412
rect 4476 124684 4740 124694
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4476 124618 4740 124628
rect 2828 124180 2884 124190
rect 2828 124086 2884 124124
rect 5136 123900 5400 123910
rect 5192 123844 5240 123900
rect 5296 123844 5344 123900
rect 5136 123834 5400 123844
rect 4476 123116 4740 123126
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4476 123050 4740 123060
rect 5136 122332 5400 122342
rect 5192 122276 5240 122332
rect 5296 122276 5344 122332
rect 5136 122266 5400 122276
rect 4476 121548 4740 121558
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4476 121482 4740 121492
rect 5136 120764 5400 120774
rect 5192 120708 5240 120764
rect 5296 120708 5344 120764
rect 5136 120698 5400 120708
rect 4476 119980 4740 119990
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4476 119914 4740 119924
rect 5136 119196 5400 119206
rect 5192 119140 5240 119196
rect 5296 119140 5344 119196
rect 5136 119130 5400 119140
rect 4476 118412 4740 118422
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4476 118346 4740 118356
rect 5136 117628 5400 117638
rect 5192 117572 5240 117628
rect 5296 117572 5344 117628
rect 5136 117562 5400 117572
rect 4476 116844 4740 116854
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4476 116778 4740 116788
rect 5136 116060 5400 116070
rect 5192 116004 5240 116060
rect 5296 116004 5344 116060
rect 5136 115994 5400 116004
rect 4476 115276 4740 115286
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4476 115210 4740 115220
rect 5136 114492 5400 114502
rect 5192 114436 5240 114492
rect 5296 114436 5344 114492
rect 5136 114426 5400 114436
rect 4476 113708 4740 113718
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4476 113642 4740 113652
rect 5136 112924 5400 112934
rect 5192 112868 5240 112924
rect 5296 112868 5344 112924
rect 5136 112858 5400 112868
rect 2828 112420 2884 112430
rect 2828 112326 2884 112364
rect 9212 112420 9268 112430
rect 4476 112140 4740 112150
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4476 112074 4740 112084
rect 5136 111356 5400 111366
rect 5192 111300 5240 111356
rect 5296 111300 5344 111356
rect 5136 111290 5400 111300
rect 4476 110572 4740 110582
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4476 110506 4740 110516
rect 5136 109788 5400 109798
rect 5192 109732 5240 109788
rect 5296 109732 5344 109788
rect 5136 109722 5400 109732
rect 4476 109004 4740 109014
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4476 108938 4740 108948
rect 5136 108220 5400 108230
rect 5192 108164 5240 108220
rect 5296 108164 5344 108220
rect 5136 108154 5400 108164
rect 4476 107436 4740 107446
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4476 107370 4740 107380
rect 5136 106652 5400 106662
rect 5192 106596 5240 106652
rect 5296 106596 5344 106652
rect 5136 106586 5400 106596
rect 4476 105868 4740 105878
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4476 105802 4740 105812
rect 5136 105084 5400 105094
rect 5192 105028 5240 105084
rect 5296 105028 5344 105084
rect 5136 105018 5400 105028
rect 4476 104300 4740 104310
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4476 104234 4740 104244
rect 5136 103516 5400 103526
rect 5192 103460 5240 103516
rect 5296 103460 5344 103516
rect 5136 103450 5400 103460
rect 4476 102732 4740 102742
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4476 102666 4740 102676
rect 5136 101948 5400 101958
rect 5192 101892 5240 101948
rect 5296 101892 5344 101948
rect 5136 101882 5400 101892
rect 7532 101668 7588 101678
rect 2492 101444 2548 101454
rect 2492 101350 2548 101388
rect 4476 101164 4740 101174
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4476 101098 4740 101108
rect 5136 100380 5400 100390
rect 5192 100324 5240 100380
rect 5296 100324 5344 100380
rect 5136 100314 5400 100324
rect 4476 99596 4740 99606
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4476 99530 4740 99540
rect 5136 98812 5400 98822
rect 5192 98756 5240 98812
rect 5296 98756 5344 98812
rect 5136 98746 5400 98756
rect 4476 98028 4740 98038
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4476 97962 4740 97972
rect 5136 97244 5400 97254
rect 5192 97188 5240 97244
rect 5296 97188 5344 97244
rect 5136 97178 5400 97188
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 5136 95676 5400 95686
rect 5192 95620 5240 95676
rect 5296 95620 5344 95676
rect 5136 95610 5400 95620
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 5136 94108 5400 94118
rect 5192 94052 5240 94108
rect 5296 94052 5344 94108
rect 5136 94042 5400 94052
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 5136 92540 5400 92550
rect 5192 92484 5240 92540
rect 5296 92484 5344 92540
rect 5136 92474 5400 92484
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 5136 90972 5400 90982
rect 5192 90916 5240 90972
rect 5296 90916 5344 90972
rect 5136 90906 5400 90916
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 2492 89570 2548 89582
rect 2492 89518 2494 89570
rect 2546 89518 2548 89570
rect 2492 89460 2548 89518
rect 2492 89394 2548 89404
rect 5136 89404 5400 89414
rect 5192 89348 5240 89404
rect 5296 89348 5344 89404
rect 5136 89338 5400 89348
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 5136 87836 5400 87846
rect 5192 87780 5240 87836
rect 5296 87780 5344 87836
rect 5136 87770 5400 87780
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 5136 86268 5400 86278
rect 5192 86212 5240 86268
rect 5296 86212 5344 86268
rect 5136 86202 5400 86212
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 5136 84700 5400 84710
rect 5192 84644 5240 84700
rect 5296 84644 5344 84700
rect 5136 84634 5400 84644
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 5136 83132 5400 83142
rect 5192 83076 5240 83132
rect 5296 83076 5344 83132
rect 5136 83066 5400 83076
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 5136 81564 5400 81574
rect 5192 81508 5240 81564
rect 5296 81508 5344 81564
rect 5136 81498 5400 81508
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 5136 79996 5400 80006
rect 5192 79940 5240 79996
rect 5296 79940 5344 79996
rect 5136 79930 5400 79940
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 2492 78596 2548 78606
rect 2492 78502 2548 78540
rect 5136 78428 5400 78438
rect 5192 78372 5240 78428
rect 5296 78372 5344 78428
rect 5136 78362 5400 78372
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 5136 76860 5400 76870
rect 5192 76804 5240 76860
rect 5296 76804 5344 76860
rect 5136 76794 5400 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 5136 75292 5400 75302
rect 5192 75236 5240 75292
rect 5296 75236 5344 75292
rect 5136 75226 5400 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 5136 73724 5400 73734
rect 5192 73668 5240 73724
rect 5296 73668 5344 73724
rect 5136 73658 5400 73668
rect 7532 73220 7588 101612
rect 7532 73154 7588 73164
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 5136 72156 5400 72166
rect 5192 72100 5240 72156
rect 5296 72100 5344 72156
rect 5136 72090 5400 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 5136 70588 5400 70598
rect 5192 70532 5240 70588
rect 5296 70532 5344 70588
rect 5136 70522 5400 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 5136 69020 5400 69030
rect 5192 68964 5240 69020
rect 5296 68964 5344 69020
rect 5136 68954 5400 68964
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 5136 67452 5400 67462
rect 5192 67396 5240 67452
rect 5296 67396 5344 67452
rect 5136 67386 5400 67396
rect 2492 66946 2548 66958
rect 2492 66894 2494 66946
rect 2546 66894 2548 66946
rect 2492 66612 2548 66894
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 2492 66546 2548 66556
rect 5136 65884 5400 65894
rect 5192 65828 5240 65884
rect 5296 65828 5344 65884
rect 5136 65818 5400 65828
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 5136 64316 5400 64326
rect 5192 64260 5240 64316
rect 5296 64260 5344 64316
rect 5136 64250 5400 64260
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 5136 62748 5400 62758
rect 5192 62692 5240 62748
rect 5296 62692 5344 62748
rect 5136 62682 5400 62692
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 5136 61180 5400 61190
rect 5192 61124 5240 61180
rect 5296 61124 5344 61180
rect 5136 61114 5400 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 5136 59612 5400 59622
rect 5192 59556 5240 59612
rect 5296 59556 5344 59612
rect 5136 59546 5400 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 5136 58044 5400 58054
rect 5192 57988 5240 58044
rect 5296 57988 5344 58044
rect 5136 57978 5400 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 5136 56476 5400 56486
rect 5192 56420 5240 56476
rect 5296 56420 5344 56476
rect 5136 56410 5400 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5136 54908 5400 54918
rect 5192 54852 5240 54908
rect 5296 54852 5344 54908
rect 5136 54842 5400 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 5136 53340 5400 53350
rect 5192 53284 5240 53340
rect 5296 53284 5344 53340
rect 5136 53274 5400 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 5136 51772 5400 51782
rect 5192 51716 5240 51772
rect 5296 51716 5344 51772
rect 5136 51706 5400 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5136 50204 5400 50214
rect 5192 50148 5240 50204
rect 5296 50148 5344 50204
rect 5136 50138 5400 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 5136 48636 5400 48646
rect 5192 48580 5240 48636
rect 5296 48580 5344 48636
rect 5136 48570 5400 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 5136 47068 5400 47078
rect 5192 47012 5240 47068
rect 5296 47012 5344 47068
rect 5136 47002 5400 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 5136 45500 5400 45510
rect 5192 45444 5240 45500
rect 5296 45444 5344 45500
rect 5136 45434 5400 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5136 43932 5400 43942
rect 5192 43876 5240 43932
rect 5296 43876 5344 43932
rect 5136 43866 5400 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5136 42364 5400 42374
rect 5192 42308 5240 42364
rect 5296 42308 5344 42364
rect 5136 42298 5400 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5136 40796 5400 40806
rect 5192 40740 5240 40796
rect 5296 40740 5344 40796
rect 5136 40730 5400 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5136 39228 5400 39238
rect 5192 39172 5240 39228
rect 5296 39172 5344 39228
rect 5136 39162 5400 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5136 37660 5400 37670
rect 5192 37604 5240 37660
rect 5296 37604 5344 37660
rect 5136 37594 5400 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 5136 36092 5400 36102
rect 5192 36036 5240 36092
rect 5296 36036 5344 36092
rect 5136 36026 5400 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5136 34524 5400 34534
rect 5192 34468 5240 34524
rect 5296 34468 5344 34524
rect 5136 34458 5400 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5136 32956 5400 32966
rect 5192 32900 5240 32956
rect 5296 32900 5344 32956
rect 5136 32890 5400 32900
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 32340 2548 32398
rect 2492 32274 2548 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5136 31388 5400 31398
rect 5192 31332 5240 31388
rect 5296 31332 5344 31388
rect 5136 31322 5400 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5136 29820 5400 29830
rect 5192 29764 5240 29820
rect 5296 29764 5344 29820
rect 5136 29754 5400 29764
rect 2380 29362 2436 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5136 28252 5400 28262
rect 5192 28196 5240 28252
rect 5296 28196 5344 28252
rect 5136 28186 5400 28196
rect 9212 27748 9268 112364
rect 9212 27682 9268 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 5136 26684 5400 26694
rect 5192 26628 5240 26684
rect 5296 26628 5344 26684
rect 5136 26618 5400 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 5136 25116 5400 25126
rect 5192 25060 5240 25116
rect 5296 25060 5344 25116
rect 5136 25050 5400 25060
rect 12572 24388 12628 146860
rect 17724 135156 17780 135166
rect 14252 78596 14308 78606
rect 14252 44324 14308 78540
rect 17612 78596 17668 78606
rect 17612 78502 17668 78540
rect 17612 77922 17668 77934
rect 17612 77870 17614 77922
rect 17666 77870 17668 77922
rect 15932 76580 15988 76590
rect 15932 55300 15988 76524
rect 17612 76580 17668 77870
rect 17612 76514 17668 76524
rect 17612 76356 17668 76366
rect 17612 76262 17668 76300
rect 17500 75684 17556 75694
rect 17500 75590 17556 75628
rect 17500 74788 17556 74798
rect 17500 74694 17556 74732
rect 17500 73220 17556 73230
rect 17500 73126 17556 73164
rect 15932 55234 15988 55244
rect 14252 44258 14308 44268
rect 17612 36260 17668 36270
rect 17612 36166 17668 36204
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 12572 24322 12628 24332
rect 12684 35588 12740 35598
rect 4476 24266 4740 24276
rect 5136 23548 5400 23558
rect 5192 23492 5240 23548
rect 5296 23492 5344 23548
rect 5136 23482 5400 23492
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5136 21980 5400 21990
rect 5192 21924 5240 21980
rect 5296 21924 5344 21980
rect 5136 21914 5400 21924
rect 2044 21810 2212 21812
rect 2044 21758 2046 21810
rect 2098 21758 2212 21810
rect 2044 21756 2212 21758
rect 2044 21746 2100 21756
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21476 1764 21534
rect 1708 20916 1764 21420
rect 2492 21476 2548 21486
rect 2492 21382 2548 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1708 20850 1764 20860
rect 5136 20412 5400 20422
rect 5192 20356 5240 20412
rect 5296 20356 5344 20412
rect 5136 20346 5400 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 5136 18844 5400 18854
rect 5192 18788 5240 18844
rect 5296 18788 5344 18844
rect 5136 18778 5400 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1708 17442 1764 17454
rect 1708 17390 1710 17442
rect 1762 17390 1764 17442
rect 1708 17108 1764 17390
rect 5136 17276 5400 17286
rect 5192 17220 5240 17276
rect 5296 17220 5344 17276
rect 5136 17210 5400 17220
rect 1708 17042 1764 17052
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5136 15708 5400 15718
rect 5192 15652 5240 15708
rect 5296 15652 5344 15708
rect 5136 15642 5400 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5136 14140 5400 14150
rect 5192 14084 5240 14140
rect 5296 14084 5344 14140
rect 5136 14074 5400 14084
rect 1708 13522 1764 13534
rect 1708 13470 1710 13522
rect 1762 13470 1764 13522
rect 1708 13300 1764 13470
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 1708 13234 1764 13244
rect 5136 12572 5400 12582
rect 5192 12516 5240 12572
rect 5296 12516 5344 12572
rect 5136 12506 5400 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5136 11004 5400 11014
rect 5192 10948 5240 11004
rect 5296 10948 5344 11004
rect 5136 10938 5400 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1708 9602 1764 9614
rect 1708 9550 1710 9602
rect 1762 9550 1764 9602
rect 1708 9492 1764 9550
rect 2044 9604 2100 9614
rect 2044 9510 2100 9548
rect 2492 9602 2548 9614
rect 2492 9550 2494 9602
rect 2546 9550 2548 9602
rect 1708 9426 1764 9436
rect 2492 9492 2548 9550
rect 12684 9604 12740 35532
rect 16940 35586 16996 35598
rect 16940 35534 16942 35586
rect 16994 35534 16996 35586
rect 16940 34692 16996 35534
rect 17612 35588 17668 35598
rect 17612 35494 17668 35532
rect 16940 34626 16996 34636
rect 17724 20468 17780 135100
rect 17724 20402 17780 20412
rect 22764 18452 22820 156268
rect 26684 156212 26740 159264
rect 34300 156660 34356 159264
rect 35856 156828 36120 156838
rect 35912 156772 35960 156828
rect 36016 156772 36064 156828
rect 35856 156762 36120 156772
rect 34524 156660 34580 156670
rect 34300 156658 34580 156660
rect 34300 156606 34526 156658
rect 34578 156606 34580 156658
rect 34300 156604 34580 156606
rect 34524 156594 34580 156604
rect 41916 156660 41972 159264
rect 41916 156434 41972 156604
rect 43708 156660 43764 156670
rect 43708 156566 43764 156604
rect 41916 156382 41918 156434
rect 41970 156382 41972 156434
rect 41916 156370 41972 156382
rect 42812 156324 42868 156334
rect 42812 156230 42868 156268
rect 26908 156212 26964 156222
rect 26684 156210 26964 156212
rect 26684 156158 26910 156210
rect 26962 156158 26964 156210
rect 26684 156156 26964 156158
rect 49532 156212 49588 159264
rect 57148 156660 57204 159264
rect 57372 156660 57428 156670
rect 57148 156658 57428 156660
rect 57148 156606 57374 156658
rect 57426 156606 57428 156658
rect 57148 156604 57428 156606
rect 57372 156594 57428 156604
rect 64764 156660 64820 159264
rect 66576 156828 66840 156838
rect 66632 156772 66680 156828
rect 66736 156772 66784 156828
rect 66576 156762 66840 156772
rect 63756 156548 63812 156558
rect 56252 156324 56308 156334
rect 49756 156212 49812 156222
rect 49532 156210 49812 156212
rect 49532 156158 49758 156210
rect 49810 156158 49812 156210
rect 49532 156156 49812 156158
rect 26908 156146 26964 156156
rect 49756 156146 49812 156156
rect 35196 156044 35460 156054
rect 35252 155988 35300 156044
rect 35356 155988 35404 156044
rect 35196 155978 35460 155988
rect 35856 155260 36120 155270
rect 35912 155204 35960 155260
rect 36016 155204 36064 155260
rect 35856 155194 36120 155204
rect 35196 154476 35460 154486
rect 35252 154420 35300 154476
rect 35356 154420 35404 154476
rect 35196 154410 35460 154420
rect 35856 153692 36120 153702
rect 35912 153636 35960 153692
rect 36016 153636 36064 153692
rect 35856 153626 36120 153636
rect 35196 152908 35460 152918
rect 35252 152852 35300 152908
rect 35356 152852 35404 152908
rect 35196 152842 35460 152852
rect 35856 152124 36120 152134
rect 35912 152068 35960 152124
rect 36016 152068 36064 152124
rect 35856 152058 36120 152068
rect 35196 151340 35460 151350
rect 35252 151284 35300 151340
rect 35356 151284 35404 151340
rect 35196 151274 35460 151284
rect 35856 150556 36120 150566
rect 35912 150500 35960 150556
rect 36016 150500 36064 150556
rect 35856 150490 36120 150500
rect 35196 149772 35460 149782
rect 35252 149716 35300 149772
rect 35356 149716 35404 149772
rect 35196 149706 35460 149716
rect 35856 148988 36120 148998
rect 35912 148932 35960 148988
rect 36016 148932 36064 148988
rect 35856 148922 36120 148932
rect 35196 148204 35460 148214
rect 35252 148148 35300 148204
rect 35356 148148 35404 148204
rect 35196 148138 35460 148148
rect 35856 147420 36120 147430
rect 35912 147364 35960 147420
rect 36016 147364 36064 147420
rect 35856 147354 36120 147364
rect 35196 146636 35460 146646
rect 35252 146580 35300 146636
rect 35356 146580 35404 146636
rect 35196 146570 35460 146580
rect 35856 145852 36120 145862
rect 35912 145796 35960 145852
rect 36016 145796 36064 145852
rect 35856 145786 36120 145796
rect 35196 145068 35460 145078
rect 35252 145012 35300 145068
rect 35356 145012 35404 145068
rect 35196 145002 35460 145012
rect 26012 124180 26068 124190
rect 26012 38052 26068 124124
rect 56252 41188 56308 156268
rect 56252 41122 56308 41132
rect 63756 41076 63812 156492
rect 64764 156434 64820 156604
rect 66556 156660 66612 156670
rect 66556 156566 66612 156604
rect 64764 156382 64766 156434
rect 64818 156382 64820 156434
rect 64764 156370 64820 156382
rect 65100 156436 65156 156446
rect 64428 156324 64484 156334
rect 64428 41300 64484 156268
rect 64428 41234 64484 41244
rect 63756 41010 63812 41020
rect 61740 38164 61796 38174
rect 26012 37986 26068 37996
rect 51436 38052 51492 38062
rect 44156 24388 44212 24398
rect 44156 21812 44212 24332
rect 51436 22372 51492 37996
rect 59052 38052 59108 38062
rect 53900 27748 53956 27758
rect 51492 22316 51604 22372
rect 51436 22306 51492 22316
rect 44156 21746 44212 21756
rect 22764 18386 22820 18396
rect 44716 21252 44772 21262
rect 35856 17276 36120 17286
rect 35912 17220 35960 17276
rect 36016 17220 36064 17276
rect 35856 17210 36120 17220
rect 44716 17106 44772 21196
rect 48300 20468 48356 20478
rect 48300 20188 48356 20412
rect 44716 17054 44718 17106
rect 44770 17054 44772 17106
rect 44716 17042 44772 17054
rect 48188 20132 48356 20188
rect 48188 17106 48244 20132
rect 48188 17054 48190 17106
rect 48242 17054 48244 17106
rect 48188 17042 48244 17054
rect 51548 17106 51604 22316
rect 53900 21812 53956 27692
rect 53900 21746 53956 21756
rect 51548 17054 51550 17106
rect 51602 17054 51604 17106
rect 51548 17042 51604 17054
rect 55132 21700 55188 21710
rect 55132 17106 55188 21644
rect 55132 17054 55134 17106
rect 55186 17054 55188 17106
rect 55132 17042 55188 17054
rect 59052 19908 59108 37996
rect 61740 22372 61796 38108
rect 61740 20188 61796 22316
rect 65100 22372 65156 156380
rect 65324 156324 65380 156334
rect 65324 156230 65380 156268
rect 72380 156212 72436 159264
rect 79996 156660 80052 159264
rect 87612 157106 87668 159264
rect 87612 157054 87614 157106
rect 87666 157054 87668 157106
rect 87612 157042 87668 157054
rect 88508 157106 88564 157118
rect 88508 157054 88510 157106
rect 88562 157054 88564 157106
rect 80220 156660 80276 156670
rect 79996 156658 80276 156660
rect 79996 156606 80222 156658
rect 80274 156606 80276 156658
rect 79996 156604 80276 156606
rect 80220 156594 80276 156604
rect 87612 156548 87668 156558
rect 87612 156454 87668 156492
rect 88508 156434 88564 157054
rect 89404 157106 89460 157118
rect 89404 157054 89406 157106
rect 89458 157054 89460 157106
rect 89404 156658 89460 157054
rect 89404 156606 89406 156658
rect 89458 156606 89460 156658
rect 89404 156594 89460 156606
rect 88508 156382 88510 156434
rect 88562 156382 88564 156434
rect 88508 156370 88564 156382
rect 72604 156212 72660 156222
rect 72380 156210 72660 156212
rect 72380 156158 72606 156210
rect 72658 156158 72660 156210
rect 72380 156156 72660 156158
rect 95228 156212 95284 159264
rect 97296 156828 97560 156838
rect 97352 156772 97400 156828
rect 97456 156772 97504 156828
rect 97296 156762 97560 156772
rect 102844 156660 102900 159264
rect 103068 156660 103124 156670
rect 102844 156658 103124 156660
rect 102844 156606 103070 156658
rect 103122 156606 103124 156658
rect 102844 156604 103124 156606
rect 103068 156594 103124 156604
rect 110460 156660 110516 159264
rect 110684 156660 110740 156670
rect 110460 156658 110740 156660
rect 110460 156606 110462 156658
rect 110514 156606 110686 156658
rect 110738 156606 110740 156658
rect 110460 156604 110740 156606
rect 110460 156594 110516 156604
rect 110684 156594 110740 156604
rect 111132 156324 111188 156334
rect 111132 156230 111188 156268
rect 95452 156212 95508 156222
rect 95228 156210 95508 156212
rect 95228 156158 95454 156210
rect 95506 156158 95508 156210
rect 95228 156156 95508 156158
rect 118076 156212 118132 159264
rect 125692 156660 125748 159264
rect 133308 157442 133364 159264
rect 133308 157390 133310 157442
rect 133362 157390 133364 157442
rect 133308 157378 133364 157390
rect 134204 157442 134260 157454
rect 134204 157390 134206 157442
rect 134258 157390 134260 157442
rect 128016 156828 128280 156838
rect 128072 156772 128120 156828
rect 128176 156772 128224 156828
rect 128016 156762 128280 156772
rect 125916 156660 125972 156670
rect 125692 156658 125972 156660
rect 125692 156606 125918 156658
rect 125970 156606 125972 156658
rect 125692 156604 125972 156606
rect 125916 156594 125972 156604
rect 134204 156660 134260 157390
rect 134204 156434 134260 156604
rect 135100 156660 135156 156670
rect 135100 156566 135156 156604
rect 134204 156382 134206 156434
rect 134258 156382 134260 156434
rect 134204 156370 134260 156382
rect 118300 156212 118356 156222
rect 118076 156210 118356 156212
rect 118076 156158 118302 156210
rect 118354 156158 118356 156210
rect 118076 156156 118356 156158
rect 72604 156146 72660 156156
rect 95452 156146 95508 156156
rect 118300 156146 118356 156156
rect 133420 156210 133476 156222
rect 133420 156158 133422 156210
rect 133474 156158 133476 156210
rect 65916 156044 66180 156054
rect 65972 155988 66020 156044
rect 66076 155988 66124 156044
rect 65916 155978 66180 155988
rect 96636 156044 96900 156054
rect 96692 155988 96740 156044
rect 96796 155988 96844 156044
rect 96636 155978 96900 155988
rect 127356 156044 127620 156054
rect 127412 155988 127460 156044
rect 127516 155988 127564 156044
rect 127356 155978 127620 155988
rect 66576 155260 66840 155270
rect 66632 155204 66680 155260
rect 66736 155204 66784 155260
rect 66576 155194 66840 155204
rect 97296 155260 97560 155270
rect 97352 155204 97400 155260
rect 97456 155204 97504 155260
rect 97296 155194 97560 155204
rect 128016 155260 128280 155270
rect 128072 155204 128120 155260
rect 128176 155204 128224 155260
rect 128016 155194 128280 155204
rect 65916 154476 66180 154486
rect 65972 154420 66020 154476
rect 66076 154420 66124 154476
rect 65916 154410 66180 154420
rect 96636 154476 96900 154486
rect 96692 154420 96740 154476
rect 96796 154420 96844 154476
rect 96636 154410 96900 154420
rect 127356 154476 127620 154486
rect 127412 154420 127460 154476
rect 127516 154420 127564 154476
rect 127356 154410 127620 154420
rect 66576 153692 66840 153702
rect 66632 153636 66680 153692
rect 66736 153636 66784 153692
rect 66576 153626 66840 153636
rect 97296 153692 97560 153702
rect 97352 153636 97400 153692
rect 97456 153636 97504 153692
rect 97296 153626 97560 153636
rect 128016 153692 128280 153702
rect 128072 153636 128120 153692
rect 128176 153636 128224 153692
rect 128016 153626 128280 153636
rect 65916 152908 66180 152918
rect 65972 152852 66020 152908
rect 66076 152852 66124 152908
rect 65916 152842 66180 152852
rect 96636 152908 96900 152918
rect 96692 152852 96740 152908
rect 96796 152852 96844 152908
rect 96636 152842 96900 152852
rect 127356 152908 127620 152918
rect 127412 152852 127460 152908
rect 127516 152852 127564 152908
rect 127356 152842 127620 152852
rect 66576 152124 66840 152134
rect 66632 152068 66680 152124
rect 66736 152068 66784 152124
rect 66576 152058 66840 152068
rect 97296 152124 97560 152134
rect 97352 152068 97400 152124
rect 97456 152068 97504 152124
rect 97296 152058 97560 152068
rect 128016 152124 128280 152134
rect 128072 152068 128120 152124
rect 128176 152068 128224 152124
rect 128016 152058 128280 152068
rect 65916 151340 66180 151350
rect 65972 151284 66020 151340
rect 66076 151284 66124 151340
rect 65916 151274 66180 151284
rect 96636 151340 96900 151350
rect 96692 151284 96740 151340
rect 96796 151284 96844 151340
rect 96636 151274 96900 151284
rect 127356 151340 127620 151350
rect 127412 151284 127460 151340
rect 127516 151284 127564 151340
rect 127356 151274 127620 151284
rect 66576 150556 66840 150566
rect 66632 150500 66680 150556
rect 66736 150500 66784 150556
rect 66576 150490 66840 150500
rect 97296 150556 97560 150566
rect 97352 150500 97400 150556
rect 97456 150500 97504 150556
rect 97296 150490 97560 150500
rect 128016 150556 128280 150566
rect 128072 150500 128120 150556
rect 128176 150500 128224 150556
rect 128016 150490 128280 150500
rect 65916 149772 66180 149782
rect 65972 149716 66020 149772
rect 66076 149716 66124 149772
rect 65916 149706 66180 149716
rect 96636 149772 96900 149782
rect 96692 149716 96740 149772
rect 96796 149716 96844 149772
rect 96636 149706 96900 149716
rect 127356 149772 127620 149782
rect 127412 149716 127460 149772
rect 127516 149716 127564 149772
rect 127356 149706 127620 149716
rect 133420 149548 133476 156158
rect 140924 156212 140980 159264
rect 148540 156660 148596 159264
rect 156156 157108 156212 159264
rect 156268 157108 156324 157118
rect 156156 157106 156324 157108
rect 156156 157054 156270 157106
rect 156322 157054 156324 157106
rect 156156 157052 156324 157054
rect 156268 157042 156324 157052
rect 157052 157106 157108 157118
rect 157052 157054 157054 157106
rect 157106 157054 157108 157106
rect 148764 156660 148820 156670
rect 148540 156658 148820 156660
rect 148540 156606 148766 156658
rect 148818 156606 148820 156658
rect 148540 156604 148820 156606
rect 148764 156594 148820 156604
rect 157052 156434 157108 157054
rect 157948 157106 158004 157118
rect 157948 157054 157950 157106
rect 158002 157054 158004 157106
rect 157948 156658 158004 157054
rect 158736 156828 159000 156838
rect 158792 156772 158840 156828
rect 158896 156772 158944 156828
rect 158736 156762 159000 156772
rect 157948 156606 157950 156658
rect 158002 156606 158004 156658
rect 157948 156594 158004 156606
rect 163772 156660 163828 159264
rect 171388 157444 171444 159264
rect 171388 157388 171892 157444
rect 163996 156660 164052 156670
rect 163772 156658 164052 156660
rect 163772 156606 163998 156658
rect 164050 156606 164052 156658
rect 163772 156604 164052 156606
rect 163996 156594 164052 156604
rect 157052 156382 157054 156434
rect 157106 156382 157108 156434
rect 157052 156370 157108 156382
rect 156380 156322 156436 156334
rect 156380 156270 156382 156322
rect 156434 156270 156436 156322
rect 141148 156212 141204 156222
rect 140924 156210 141204 156212
rect 140924 156158 141150 156210
rect 141202 156158 141204 156210
rect 140924 156156 141204 156158
rect 141148 156146 141204 156156
rect 132972 149492 133476 149548
rect 66576 148988 66840 148998
rect 66632 148932 66680 148988
rect 66736 148932 66784 148988
rect 66576 148922 66840 148932
rect 97296 148988 97560 148998
rect 97352 148932 97400 148988
rect 97456 148932 97504 148988
rect 97296 148922 97560 148932
rect 128016 148988 128280 148998
rect 128072 148932 128120 148988
rect 128176 148932 128224 148988
rect 128016 148922 128280 148932
rect 65916 148204 66180 148214
rect 65972 148148 66020 148204
rect 66076 148148 66124 148204
rect 65916 148138 66180 148148
rect 96636 148204 96900 148214
rect 96692 148148 96740 148204
rect 96796 148148 96844 148204
rect 96636 148138 96900 148148
rect 127356 148204 127620 148214
rect 127412 148148 127460 148204
rect 127516 148148 127564 148204
rect 127356 148138 127620 148148
rect 66576 147420 66840 147430
rect 66632 147364 66680 147420
rect 66736 147364 66784 147420
rect 66576 147354 66840 147364
rect 97296 147420 97560 147430
rect 97352 147364 97400 147420
rect 97456 147364 97504 147420
rect 97296 147354 97560 147364
rect 128016 147420 128280 147430
rect 128072 147364 128120 147420
rect 128176 147364 128224 147420
rect 128016 147354 128280 147364
rect 65916 146636 66180 146646
rect 65972 146580 66020 146636
rect 66076 146580 66124 146636
rect 65916 146570 66180 146580
rect 96636 146636 96900 146646
rect 96692 146580 96740 146636
rect 96796 146580 96844 146636
rect 96636 146570 96900 146580
rect 127356 146636 127620 146646
rect 127412 146580 127460 146636
rect 127516 146580 127564 146636
rect 127356 146570 127620 146580
rect 66576 145852 66840 145862
rect 66632 145796 66680 145852
rect 66736 145796 66784 145852
rect 66576 145786 66840 145796
rect 97296 145852 97560 145862
rect 97352 145796 97400 145852
rect 97456 145796 97504 145852
rect 97296 145786 97560 145796
rect 128016 145852 128280 145862
rect 128072 145796 128120 145852
rect 128176 145796 128224 145852
rect 128016 145786 128280 145796
rect 65916 145068 66180 145078
rect 65972 145012 66020 145068
rect 66076 145012 66124 145068
rect 65916 145002 66180 145012
rect 96636 145068 96900 145078
rect 96692 145012 96740 145068
rect 96796 145012 96844 145068
rect 96636 145002 96900 145012
rect 127356 145068 127620 145078
rect 127412 145012 127460 145068
rect 127516 145012 127564 145068
rect 127356 145002 127620 145012
rect 132972 47012 133028 149492
rect 132972 46946 133028 46956
rect 156380 47012 156436 156270
rect 158076 156044 158340 156054
rect 158132 155988 158180 156044
rect 158236 155988 158284 156044
rect 158076 155978 158340 155988
rect 171836 155874 171892 157388
rect 186620 156660 186676 159264
rect 189456 156828 189720 156838
rect 189512 156772 189560 156828
rect 189616 156772 189664 156828
rect 189456 156762 189720 156772
rect 186844 156660 186900 156670
rect 186620 156658 186900 156660
rect 186620 156606 186846 156658
rect 186898 156606 186900 156658
rect 186620 156604 186900 156606
rect 186844 156594 186900 156604
rect 188796 156044 189060 156054
rect 188852 155988 188900 156044
rect 188956 155988 189004 156044
rect 188796 155978 189060 155988
rect 171836 155822 171838 155874
rect 171890 155822 171892 155874
rect 171836 155810 171892 155822
rect 194236 155876 194292 159264
rect 194236 155810 194292 155820
rect 194908 155876 194964 155886
rect 194908 155762 194964 155820
rect 194908 155710 194910 155762
rect 194962 155710 194964 155762
rect 194908 155698 194964 155710
rect 174188 155650 174244 155662
rect 174188 155598 174190 155650
rect 174242 155598 174244 155650
rect 174188 155428 174244 155598
rect 196588 155650 196644 155662
rect 196588 155598 196590 155650
rect 196642 155598 196644 155650
rect 174636 155428 174692 155438
rect 174188 155426 174692 155428
rect 174188 155374 174638 155426
rect 174690 155374 174692 155426
rect 174188 155372 174692 155374
rect 158736 155260 159000 155270
rect 158792 155204 158840 155260
rect 158896 155204 158944 155260
rect 158736 155194 159000 155204
rect 158076 154476 158340 154486
rect 158132 154420 158180 154476
rect 158236 154420 158284 154476
rect 158076 154410 158340 154420
rect 158736 153692 159000 153702
rect 158792 153636 158840 153692
rect 158896 153636 158944 153692
rect 158736 153626 159000 153636
rect 158076 152908 158340 152918
rect 158132 152852 158180 152908
rect 158236 152852 158284 152908
rect 158076 152842 158340 152852
rect 158736 152124 159000 152134
rect 158792 152068 158840 152124
rect 158896 152068 158944 152124
rect 158736 152058 159000 152068
rect 158076 151340 158340 151350
rect 158132 151284 158180 151340
rect 158236 151284 158284 151340
rect 158076 151274 158340 151284
rect 158736 150556 159000 150566
rect 158792 150500 158840 150556
rect 158896 150500 158944 150556
rect 158736 150490 159000 150500
rect 158076 149772 158340 149782
rect 158132 149716 158180 149772
rect 158236 149716 158284 149772
rect 158076 149706 158340 149716
rect 174636 149548 174692 155372
rect 196588 155428 196644 155598
rect 197484 155428 197540 155438
rect 196588 155426 197540 155428
rect 196588 155374 197486 155426
rect 197538 155374 197540 155426
rect 196588 155372 197540 155374
rect 189456 155260 189720 155270
rect 189512 155204 189560 155260
rect 189616 155204 189664 155260
rect 189456 155194 189720 155204
rect 188796 154476 189060 154486
rect 188852 154420 188900 154476
rect 188956 154420 189004 154476
rect 188796 154410 189060 154420
rect 189456 153692 189720 153702
rect 189512 153636 189560 153692
rect 189616 153636 189664 153692
rect 189456 153626 189720 153636
rect 188796 152908 189060 152918
rect 188852 152852 188900 152908
rect 188956 152852 189004 152908
rect 188796 152842 189060 152852
rect 189456 152124 189720 152134
rect 189512 152068 189560 152124
rect 189616 152068 189664 152124
rect 189456 152058 189720 152068
rect 188796 151340 189060 151350
rect 188852 151284 188900 151340
rect 188956 151284 189004 151340
rect 188796 151274 189060 151284
rect 189456 150556 189720 150566
rect 189512 150500 189560 150556
rect 189616 150500 189664 150556
rect 189456 150490 189720 150500
rect 188796 149772 189060 149782
rect 188852 149716 188900 149772
rect 188956 149716 189004 149772
rect 188796 149706 189060 149716
rect 174412 149492 174692 149548
rect 158736 148988 159000 148998
rect 158792 148932 158840 148988
rect 158896 148932 158944 148988
rect 158736 148922 159000 148932
rect 158076 148204 158340 148214
rect 158132 148148 158180 148204
rect 158236 148148 158284 148204
rect 158076 148138 158340 148148
rect 158736 147420 159000 147430
rect 158792 147364 158840 147420
rect 158896 147364 158944 147420
rect 158736 147354 159000 147364
rect 158076 146636 158340 146646
rect 158132 146580 158180 146636
rect 158236 146580 158284 146636
rect 158076 146570 158340 146580
rect 158736 145852 159000 145862
rect 158792 145796 158840 145852
rect 158896 145796 158944 145852
rect 158736 145786 159000 145796
rect 158076 145068 158340 145078
rect 158132 145012 158180 145068
rect 158236 145012 158284 145068
rect 158076 145002 158340 145012
rect 156380 46946 156436 46956
rect 173964 47234 174020 47246
rect 173964 47182 173966 47234
rect 174018 47182 174020 47234
rect 132972 45780 133028 45790
rect 71932 41300 71988 41310
rect 67676 41076 67732 41086
rect 65156 22316 65492 22372
rect 65100 22306 65156 22316
rect 61740 20132 62020 20188
rect 59052 17106 59108 19852
rect 59052 17054 59054 17106
rect 59106 17054 59108 17106
rect 59052 17042 59108 17054
rect 61964 17106 62020 20132
rect 61964 17054 61966 17106
rect 62018 17054 62020 17106
rect 61964 17042 62020 17054
rect 65436 17106 65492 22316
rect 67676 21812 67732 41020
rect 71932 22372 71988 41244
rect 75516 41188 75572 41198
rect 71988 22316 72100 22372
rect 71932 22306 71988 22316
rect 67676 21746 67732 21756
rect 68796 21812 68852 21822
rect 67788 20468 67844 20478
rect 67788 20188 67844 20412
rect 67788 20132 67956 20188
rect 66576 17276 66840 17286
rect 66632 17220 66680 17276
rect 66736 17220 66784 17276
rect 66576 17210 66840 17220
rect 65436 17054 65438 17106
rect 65490 17054 65492 17106
rect 65436 17042 65492 17054
rect 67900 16882 67956 20132
rect 68796 17106 68852 21756
rect 68796 17054 68798 17106
rect 68850 17054 68852 17106
rect 68796 17042 68852 17054
rect 72044 17108 72100 22316
rect 75516 21812 75572 41132
rect 85148 40964 85204 40974
rect 85148 31892 85204 40908
rect 132972 38164 133028 45724
rect 132972 38098 133028 38108
rect 156380 45780 156436 45790
rect 156380 38052 156436 45724
rect 173964 44324 174020 47182
rect 174412 47234 174468 149492
rect 189456 148988 189720 148998
rect 189512 148932 189560 148988
rect 189616 148932 189664 148988
rect 189456 148922 189720 148932
rect 188796 148204 189060 148214
rect 188852 148148 188900 148204
rect 188956 148148 189004 148204
rect 188796 148138 189060 148148
rect 189456 147420 189720 147430
rect 189512 147364 189560 147420
rect 189616 147364 189664 147420
rect 189456 147354 189720 147364
rect 188796 146636 189060 146646
rect 188852 146580 188900 146636
rect 188956 146580 189004 146636
rect 188796 146570 189060 146580
rect 189456 145852 189720 145862
rect 189512 145796 189560 145852
rect 189616 145796 189664 145852
rect 189456 145786 189720 145796
rect 188796 145068 189060 145078
rect 188852 145012 188900 145068
rect 188956 145012 189004 145068
rect 188796 145002 189060 145012
rect 189456 144284 189720 144294
rect 189512 144228 189560 144284
rect 189616 144228 189664 144284
rect 189456 144218 189720 144228
rect 188796 143500 189060 143510
rect 188852 143444 188900 143500
rect 188956 143444 189004 143500
rect 188796 143434 189060 143444
rect 189456 142716 189720 142726
rect 189512 142660 189560 142716
rect 189616 142660 189664 142716
rect 189456 142650 189720 142660
rect 188796 141932 189060 141942
rect 188852 141876 188900 141932
rect 188956 141876 189004 141932
rect 188796 141866 189060 141876
rect 189456 141148 189720 141158
rect 189512 141092 189560 141148
rect 189616 141092 189664 141148
rect 189456 141082 189720 141092
rect 188796 140364 189060 140374
rect 188852 140308 188900 140364
rect 188956 140308 189004 140364
rect 188796 140298 189060 140308
rect 189456 139580 189720 139590
rect 189512 139524 189560 139580
rect 189616 139524 189664 139580
rect 189456 139514 189720 139524
rect 188796 138796 189060 138806
rect 188852 138740 188900 138796
rect 188956 138740 189004 138796
rect 188796 138730 189060 138740
rect 189456 138012 189720 138022
rect 189512 137956 189560 138012
rect 189616 137956 189664 138012
rect 189456 137946 189720 137956
rect 188796 137228 189060 137238
rect 188852 137172 188900 137228
rect 188956 137172 189004 137228
rect 188796 137162 189060 137172
rect 189456 136444 189720 136454
rect 189512 136388 189560 136444
rect 189616 136388 189664 136444
rect 189456 136378 189720 136388
rect 188796 135660 189060 135670
rect 188852 135604 188900 135660
rect 188956 135604 189004 135660
rect 188796 135594 189060 135604
rect 189456 134876 189720 134886
rect 189512 134820 189560 134876
rect 189616 134820 189664 134876
rect 189456 134810 189720 134820
rect 188796 134092 189060 134102
rect 188852 134036 188900 134092
rect 188956 134036 189004 134092
rect 188796 134026 189060 134036
rect 189456 133308 189720 133318
rect 189512 133252 189560 133308
rect 189616 133252 189664 133308
rect 189456 133242 189720 133252
rect 188796 132524 189060 132534
rect 188852 132468 188900 132524
rect 188956 132468 189004 132524
rect 188796 132458 189060 132468
rect 189456 131740 189720 131750
rect 189512 131684 189560 131740
rect 189616 131684 189664 131740
rect 189456 131674 189720 131684
rect 188796 130956 189060 130966
rect 188852 130900 188900 130956
rect 188956 130900 189004 130956
rect 188796 130890 189060 130900
rect 189456 130172 189720 130182
rect 189512 130116 189560 130172
rect 189616 130116 189664 130172
rect 189456 130106 189720 130116
rect 188796 129388 189060 129398
rect 188852 129332 188900 129388
rect 188956 129332 189004 129388
rect 188796 129322 189060 129332
rect 189456 128604 189720 128614
rect 189512 128548 189560 128604
rect 189616 128548 189664 128604
rect 189456 128538 189720 128548
rect 188796 127820 189060 127830
rect 188852 127764 188900 127820
rect 188956 127764 189004 127820
rect 188796 127754 189060 127764
rect 189456 127036 189720 127046
rect 189512 126980 189560 127036
rect 189616 126980 189664 127036
rect 189456 126970 189720 126980
rect 188796 126252 189060 126262
rect 188852 126196 188900 126252
rect 188956 126196 189004 126252
rect 188796 126186 189060 126196
rect 189456 125468 189720 125478
rect 189512 125412 189560 125468
rect 189616 125412 189664 125468
rect 189456 125402 189720 125412
rect 188796 124684 189060 124694
rect 188852 124628 188900 124684
rect 188956 124628 189004 124684
rect 188796 124618 189060 124628
rect 189456 123900 189720 123910
rect 189512 123844 189560 123900
rect 189616 123844 189664 123900
rect 189456 123834 189720 123844
rect 188796 123116 189060 123126
rect 188852 123060 188900 123116
rect 188956 123060 189004 123116
rect 188796 123050 189060 123060
rect 189456 122332 189720 122342
rect 189512 122276 189560 122332
rect 189616 122276 189664 122332
rect 189456 122266 189720 122276
rect 188796 121548 189060 121558
rect 188852 121492 188900 121548
rect 188956 121492 189004 121548
rect 188796 121482 189060 121492
rect 189456 120764 189720 120774
rect 189512 120708 189560 120764
rect 189616 120708 189664 120764
rect 189456 120698 189720 120708
rect 188796 119980 189060 119990
rect 188852 119924 188900 119980
rect 188956 119924 189004 119980
rect 188796 119914 189060 119924
rect 189456 119196 189720 119206
rect 189512 119140 189560 119196
rect 189616 119140 189664 119196
rect 189456 119130 189720 119140
rect 188796 118412 189060 118422
rect 188852 118356 188900 118412
rect 188956 118356 189004 118412
rect 188796 118346 189060 118356
rect 189456 117628 189720 117638
rect 189512 117572 189560 117628
rect 189616 117572 189664 117628
rect 189456 117562 189720 117572
rect 188796 116844 189060 116854
rect 188852 116788 188900 116844
rect 188956 116788 189004 116844
rect 188796 116778 189060 116788
rect 189456 116060 189720 116070
rect 189512 116004 189560 116060
rect 189616 116004 189664 116060
rect 189456 115994 189720 116004
rect 188796 115276 189060 115286
rect 188852 115220 188900 115276
rect 188956 115220 189004 115276
rect 188796 115210 189060 115220
rect 189456 114492 189720 114502
rect 189512 114436 189560 114492
rect 189616 114436 189664 114492
rect 189456 114426 189720 114436
rect 188796 113708 189060 113718
rect 188852 113652 188900 113708
rect 188956 113652 189004 113708
rect 188796 113642 189060 113652
rect 189456 112924 189720 112934
rect 189512 112868 189560 112924
rect 189616 112868 189664 112924
rect 189456 112858 189720 112868
rect 188796 112140 189060 112150
rect 188852 112084 188900 112140
rect 188956 112084 189004 112140
rect 188796 112074 189060 112084
rect 189456 111356 189720 111366
rect 189512 111300 189560 111356
rect 189616 111300 189664 111356
rect 189456 111290 189720 111300
rect 188796 110572 189060 110582
rect 188852 110516 188900 110572
rect 188956 110516 189004 110572
rect 188796 110506 189060 110516
rect 189456 109788 189720 109798
rect 189512 109732 189560 109788
rect 189616 109732 189664 109788
rect 189456 109722 189720 109732
rect 188796 109004 189060 109014
rect 188852 108948 188900 109004
rect 188956 108948 189004 109004
rect 188796 108938 189060 108948
rect 189456 108220 189720 108230
rect 189512 108164 189560 108220
rect 189616 108164 189664 108220
rect 189456 108154 189720 108164
rect 188796 107436 189060 107446
rect 188852 107380 188900 107436
rect 188956 107380 189004 107436
rect 188796 107370 189060 107380
rect 189456 106652 189720 106662
rect 189512 106596 189560 106652
rect 189616 106596 189664 106652
rect 189456 106586 189720 106596
rect 188796 105868 189060 105878
rect 188852 105812 188900 105868
rect 188956 105812 189004 105868
rect 188796 105802 189060 105812
rect 189456 105084 189720 105094
rect 189512 105028 189560 105084
rect 189616 105028 189664 105084
rect 189456 105018 189720 105028
rect 188796 104300 189060 104310
rect 188852 104244 188900 104300
rect 188956 104244 189004 104300
rect 188796 104234 189060 104244
rect 189456 103516 189720 103526
rect 189512 103460 189560 103516
rect 189616 103460 189664 103516
rect 189456 103450 189720 103460
rect 188796 102732 189060 102742
rect 188852 102676 188900 102732
rect 188956 102676 189004 102732
rect 188796 102666 189060 102676
rect 189456 101948 189720 101958
rect 189512 101892 189560 101948
rect 189616 101892 189664 101948
rect 189456 101882 189720 101892
rect 188796 101164 189060 101174
rect 188852 101108 188900 101164
rect 188956 101108 189004 101164
rect 188796 101098 189060 101108
rect 189456 100380 189720 100390
rect 189512 100324 189560 100380
rect 189616 100324 189664 100380
rect 189456 100314 189720 100324
rect 188796 99596 189060 99606
rect 188852 99540 188900 99596
rect 188956 99540 189004 99596
rect 188796 99530 189060 99540
rect 189456 98812 189720 98822
rect 189512 98756 189560 98812
rect 189616 98756 189664 98812
rect 189456 98746 189720 98756
rect 188796 98028 189060 98038
rect 188852 97972 188900 98028
rect 188956 97972 189004 98028
rect 188796 97962 189060 97972
rect 189456 97244 189720 97254
rect 189512 97188 189560 97244
rect 189616 97188 189664 97244
rect 189456 97178 189720 97188
rect 188796 96460 189060 96470
rect 188852 96404 188900 96460
rect 188956 96404 189004 96460
rect 188796 96394 189060 96404
rect 189456 95676 189720 95686
rect 189512 95620 189560 95676
rect 189616 95620 189664 95676
rect 189456 95610 189720 95620
rect 188796 94892 189060 94902
rect 188852 94836 188900 94892
rect 188956 94836 189004 94892
rect 188796 94826 189060 94836
rect 189456 94108 189720 94118
rect 189512 94052 189560 94108
rect 189616 94052 189664 94108
rect 189456 94042 189720 94052
rect 190652 93716 190708 93726
rect 188796 93324 189060 93334
rect 188852 93268 188900 93324
rect 188956 93268 189004 93324
rect 188796 93258 189060 93268
rect 189456 92540 189720 92550
rect 189512 92484 189560 92540
rect 189616 92484 189664 92540
rect 189456 92474 189720 92484
rect 188796 91756 189060 91766
rect 188852 91700 188900 91756
rect 188956 91700 189004 91756
rect 188796 91690 189060 91700
rect 189456 90972 189720 90982
rect 189512 90916 189560 90972
rect 189616 90916 189664 90972
rect 189456 90906 189720 90916
rect 188796 90188 189060 90198
rect 188852 90132 188900 90188
rect 188956 90132 189004 90188
rect 188796 90122 189060 90132
rect 189456 89404 189720 89414
rect 189512 89348 189560 89404
rect 189616 89348 189664 89404
rect 189456 89338 189720 89348
rect 188796 88620 189060 88630
rect 188852 88564 188900 88620
rect 188956 88564 189004 88620
rect 188796 88554 189060 88564
rect 189456 87836 189720 87846
rect 189512 87780 189560 87836
rect 189616 87780 189664 87836
rect 189456 87770 189720 87780
rect 188796 87052 189060 87062
rect 188852 86996 188900 87052
rect 188956 86996 189004 87052
rect 188796 86986 189060 86996
rect 189456 86268 189720 86278
rect 189512 86212 189560 86268
rect 189616 86212 189664 86268
rect 189456 86202 189720 86212
rect 188796 85484 189060 85494
rect 188852 85428 188900 85484
rect 188956 85428 189004 85484
rect 188796 85418 189060 85428
rect 189456 84700 189720 84710
rect 189512 84644 189560 84700
rect 189616 84644 189664 84700
rect 189456 84634 189720 84644
rect 188796 83916 189060 83926
rect 188852 83860 188900 83916
rect 188956 83860 189004 83916
rect 188796 83850 189060 83860
rect 189456 83132 189720 83142
rect 189512 83076 189560 83132
rect 189616 83076 189664 83132
rect 189456 83066 189720 83076
rect 188796 82348 189060 82358
rect 188852 82292 188900 82348
rect 188956 82292 189004 82348
rect 188796 82282 189060 82292
rect 189456 81564 189720 81574
rect 189512 81508 189560 81564
rect 189616 81508 189664 81564
rect 189456 81498 189720 81508
rect 188796 80780 189060 80790
rect 188852 80724 188900 80780
rect 188956 80724 189004 80780
rect 188796 80714 189060 80724
rect 189456 79996 189720 80006
rect 189512 79940 189560 79996
rect 189616 79940 189664 79996
rect 189456 79930 189720 79940
rect 188796 79212 189060 79222
rect 188852 79156 188900 79212
rect 188956 79156 189004 79212
rect 188796 79146 189060 79156
rect 189456 78428 189720 78438
rect 189512 78372 189560 78428
rect 189616 78372 189664 78428
rect 189456 78362 189720 78372
rect 188796 77644 189060 77654
rect 188852 77588 188900 77644
rect 188956 77588 189004 77644
rect 188796 77578 189060 77588
rect 189456 76860 189720 76870
rect 189512 76804 189560 76860
rect 189616 76804 189664 76860
rect 189456 76794 189720 76804
rect 188796 76076 189060 76086
rect 188852 76020 188900 76076
rect 188956 76020 189004 76076
rect 188796 76010 189060 76020
rect 189456 75292 189720 75302
rect 189512 75236 189560 75292
rect 189616 75236 189664 75292
rect 189456 75226 189720 75236
rect 188796 74508 189060 74518
rect 188852 74452 188900 74508
rect 188956 74452 189004 74508
rect 188796 74442 189060 74452
rect 189456 73724 189720 73734
rect 189512 73668 189560 73724
rect 189616 73668 189664 73724
rect 189456 73658 189720 73668
rect 188796 72940 189060 72950
rect 188852 72884 188900 72940
rect 188956 72884 189004 72940
rect 188796 72874 189060 72884
rect 189456 72156 189720 72166
rect 189512 72100 189560 72156
rect 189616 72100 189664 72156
rect 189456 72090 189720 72100
rect 188796 71372 189060 71382
rect 188852 71316 188900 71372
rect 188956 71316 189004 71372
rect 188796 71306 189060 71316
rect 189456 70588 189720 70598
rect 189512 70532 189560 70588
rect 189616 70532 189664 70588
rect 189456 70522 189720 70532
rect 188796 69804 189060 69814
rect 188852 69748 188900 69804
rect 188956 69748 189004 69804
rect 188796 69738 189060 69748
rect 189456 69020 189720 69030
rect 189512 68964 189560 69020
rect 189616 68964 189664 69020
rect 189456 68954 189720 68964
rect 188796 68236 189060 68246
rect 188852 68180 188900 68236
rect 188956 68180 189004 68236
rect 188796 68170 189060 68180
rect 189456 67452 189720 67462
rect 189512 67396 189560 67452
rect 189616 67396 189664 67452
rect 189456 67386 189720 67396
rect 174412 47182 174414 47234
rect 174466 47182 174468 47234
rect 174412 47170 174468 47182
rect 187292 67060 187348 67070
rect 173964 44268 174132 44324
rect 174076 43876 174132 44268
rect 173964 43820 174132 43876
rect 173964 38724 174020 43820
rect 173964 38658 174020 38668
rect 156380 37986 156436 37996
rect 85148 31826 85204 31836
rect 72156 17108 72212 17118
rect 72044 17106 72212 17108
rect 72044 17054 72158 17106
rect 72210 17054 72212 17106
rect 72044 17052 72212 17054
rect 72156 17042 72212 17052
rect 75516 17106 75572 21756
rect 75628 29428 75684 29438
rect 75628 20468 75684 29372
rect 154588 29428 154644 29438
rect 149548 26180 149604 26190
rect 78876 25508 78932 25518
rect 78876 22708 78932 25452
rect 149548 22932 149604 26124
rect 149548 22866 149604 22876
rect 78876 22642 78932 22652
rect 97132 22708 97188 22718
rect 82908 21252 82964 21262
rect 75628 20402 75684 20412
rect 82460 20468 82516 20478
rect 82460 20188 82516 20412
rect 82348 20132 82516 20188
rect 75516 17054 75518 17106
rect 75570 17054 75572 17106
rect 75516 17042 75572 17054
rect 78988 17108 79044 17118
rect 78988 17014 79044 17052
rect 82348 17106 82404 20132
rect 82348 17054 82350 17106
rect 82402 17054 82404 17106
rect 82348 17042 82404 17054
rect 82908 17106 82964 21196
rect 82908 17054 82910 17106
rect 82962 17054 82964 17106
rect 82908 17042 82964 17054
rect 97132 17106 97188 22652
rect 140028 22708 140084 22718
rect 111244 21140 111300 21150
rect 97296 17276 97560 17286
rect 97352 17220 97400 17276
rect 97456 17220 97504 17276
rect 97296 17210 97560 17220
rect 97132 17054 97134 17106
rect 97186 17054 97188 17106
rect 97132 17042 97188 17054
rect 111244 17106 111300 21084
rect 128016 17276 128280 17286
rect 128072 17220 128120 17276
rect 128176 17220 128224 17276
rect 128016 17210 128280 17220
rect 111244 17054 111246 17106
rect 111298 17054 111300 17106
rect 111244 17042 111300 17054
rect 140028 17106 140084 22652
rect 154588 20468 154644 29372
rect 187292 25620 187348 67004
rect 188796 66668 189060 66678
rect 188852 66612 188900 66668
rect 188956 66612 189004 66668
rect 188796 66602 189060 66612
rect 189456 65884 189720 65894
rect 189512 65828 189560 65884
rect 189616 65828 189664 65884
rect 189456 65818 189720 65828
rect 188796 65100 189060 65110
rect 188852 65044 188900 65100
rect 188956 65044 189004 65100
rect 188796 65034 189060 65044
rect 189456 64316 189720 64326
rect 189512 64260 189560 64316
rect 189616 64260 189664 64316
rect 189456 64250 189720 64260
rect 188796 63532 189060 63542
rect 188852 63476 188900 63532
rect 188956 63476 189004 63532
rect 188796 63466 189060 63476
rect 189456 62748 189720 62758
rect 189512 62692 189560 62748
rect 189616 62692 189664 62748
rect 189456 62682 189720 62692
rect 188796 61964 189060 61974
rect 188852 61908 188900 61964
rect 188956 61908 189004 61964
rect 188796 61898 189060 61908
rect 189456 61180 189720 61190
rect 189512 61124 189560 61180
rect 189616 61124 189664 61180
rect 189456 61114 189720 61124
rect 188796 60396 189060 60406
rect 188852 60340 188900 60396
rect 188956 60340 189004 60396
rect 188796 60330 189060 60340
rect 189456 59612 189720 59622
rect 189512 59556 189560 59612
rect 189616 59556 189664 59612
rect 189456 59546 189720 59556
rect 188796 58828 189060 58838
rect 188852 58772 188900 58828
rect 188956 58772 189004 58828
rect 188796 58762 189060 58772
rect 189456 58044 189720 58054
rect 189512 57988 189560 58044
rect 189616 57988 189664 58044
rect 189456 57978 189720 57988
rect 188796 57260 189060 57270
rect 188852 57204 188900 57260
rect 188956 57204 189004 57260
rect 188796 57194 189060 57204
rect 189456 56476 189720 56486
rect 189512 56420 189560 56476
rect 189616 56420 189664 56476
rect 189456 56410 189720 56420
rect 188796 55692 189060 55702
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 188796 55626 189060 55636
rect 189456 54908 189720 54918
rect 189512 54852 189560 54908
rect 189616 54852 189664 54908
rect 189456 54842 189720 54852
rect 188796 54124 189060 54134
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 188796 54058 189060 54068
rect 189456 53340 189720 53350
rect 189512 53284 189560 53340
rect 189616 53284 189664 53340
rect 189456 53274 189720 53284
rect 188796 52556 189060 52566
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 188796 52490 189060 52500
rect 189456 51772 189720 51782
rect 189512 51716 189560 51772
rect 189616 51716 189664 51772
rect 189456 51706 189720 51716
rect 188796 50988 189060 50998
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 188796 50922 189060 50932
rect 189456 50204 189720 50214
rect 189512 50148 189560 50204
rect 189616 50148 189664 50204
rect 189456 50138 189720 50148
rect 188796 49420 189060 49430
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 188796 49354 189060 49364
rect 189456 48636 189720 48646
rect 189512 48580 189560 48636
rect 189616 48580 189664 48636
rect 189456 48570 189720 48580
rect 188796 47852 189060 47862
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 188796 47786 189060 47796
rect 189456 47068 189720 47078
rect 189512 47012 189560 47068
rect 189616 47012 189664 47068
rect 189456 47002 189720 47012
rect 188796 46284 189060 46294
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 188796 46218 189060 46228
rect 189456 45500 189720 45510
rect 189512 45444 189560 45500
rect 189616 45444 189664 45500
rect 189456 45434 189720 45444
rect 188796 44716 189060 44726
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 188796 44650 189060 44660
rect 189456 43932 189720 43942
rect 189512 43876 189560 43932
rect 189616 43876 189664 43932
rect 189456 43866 189720 43876
rect 188796 43148 189060 43158
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 188796 43082 189060 43092
rect 189456 42364 189720 42374
rect 189512 42308 189560 42364
rect 189616 42308 189664 42364
rect 189456 42298 189720 42308
rect 188796 41580 189060 41590
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 188796 41514 189060 41524
rect 189456 40796 189720 40806
rect 189512 40740 189560 40796
rect 189616 40740 189664 40796
rect 189456 40730 189720 40740
rect 188796 40012 189060 40022
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 188796 39946 189060 39956
rect 189456 39228 189720 39238
rect 189512 39172 189560 39228
rect 189616 39172 189664 39228
rect 189456 39162 189720 39172
rect 188748 38724 188804 38734
rect 188748 38630 188804 38668
rect 188796 38444 189060 38454
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 188796 38378 189060 38388
rect 189456 37660 189720 37670
rect 189512 37604 189560 37660
rect 189616 37604 189664 37660
rect 189456 37594 189720 37604
rect 188796 36876 189060 36886
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 188796 36810 189060 36820
rect 189456 36092 189720 36102
rect 189512 36036 189560 36092
rect 189616 36036 189664 36092
rect 189456 36026 189720 36036
rect 188796 35308 189060 35318
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 188796 35242 189060 35252
rect 189456 34524 189720 34534
rect 189512 34468 189560 34524
rect 189616 34468 189664 34524
rect 189456 34458 189720 34468
rect 188796 33740 189060 33750
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 188796 33674 189060 33684
rect 189456 32956 189720 32966
rect 189512 32900 189560 32956
rect 189616 32900 189664 32956
rect 189456 32890 189720 32900
rect 188796 32172 189060 32182
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 188796 32106 189060 32116
rect 189456 31388 189720 31398
rect 189512 31332 189560 31388
rect 189616 31332 189664 31388
rect 189456 31322 189720 31332
rect 188796 30604 189060 30614
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 188796 30538 189060 30548
rect 189456 29820 189720 29830
rect 189512 29764 189560 29820
rect 189616 29764 189664 29820
rect 189456 29754 189720 29764
rect 188796 29036 189060 29046
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 188796 28970 189060 28980
rect 189456 28252 189720 28262
rect 189512 28196 189560 28252
rect 189616 28196 189664 28252
rect 189456 28186 189720 28196
rect 188796 27468 189060 27478
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 188796 27402 189060 27412
rect 189456 26684 189720 26694
rect 189512 26628 189560 26684
rect 189616 26628 189664 26684
rect 189456 26618 189720 26628
rect 188796 25900 189060 25910
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 188796 25834 189060 25844
rect 187292 25554 187348 25564
rect 190652 25396 190708 93660
rect 196588 29428 196644 155372
rect 197484 155362 197540 155372
rect 204316 154978 204372 154990
rect 204316 154926 204318 154978
rect 204370 154926 204372 154978
rect 204316 154196 204372 154926
rect 204316 154130 204372 154140
rect 204092 146354 204148 146366
rect 204092 146302 204094 146354
rect 204146 146302 204148 146354
rect 196588 29362 196644 29372
rect 201068 146244 201124 146254
rect 201068 27860 201124 146188
rect 201740 146244 201796 146254
rect 201740 146150 201796 146188
rect 204092 145460 204148 146302
rect 204092 145394 204148 145404
rect 203756 128322 203812 128334
rect 203756 128270 203758 128322
rect 203810 128270 203812 128322
rect 203756 127988 203812 128270
rect 203756 127922 203812 127932
rect 204092 119698 204148 119710
rect 204092 119646 204094 119698
rect 204146 119646 204148 119698
rect 202188 119586 202244 119598
rect 202188 119534 202190 119586
rect 202242 119534 202244 119586
rect 202188 118692 202244 119534
rect 204092 119364 204148 119646
rect 204092 119298 204148 119308
rect 202188 114268 202244 118636
rect 203756 118692 203812 118702
rect 203756 118598 203812 118636
rect 202188 114212 202468 114268
rect 201180 93716 201236 93726
rect 201180 93622 201236 93660
rect 201180 67060 201236 67070
rect 201180 66966 201236 67004
rect 201740 41186 201796 41198
rect 201740 41134 201742 41186
rect 201794 41134 201796 41186
rect 201404 40964 201460 40974
rect 201740 40964 201796 41134
rect 201460 40908 201796 40964
rect 201404 40870 201460 40908
rect 201068 27794 201124 27804
rect 202412 27748 202468 114212
rect 204316 102114 204372 102126
rect 204316 102062 204318 102114
rect 204370 102062 204372 102114
rect 204316 101780 204372 102062
rect 204316 101714 204372 101724
rect 203980 93716 204036 93726
rect 203196 93602 203252 93614
rect 203196 93550 203198 93602
rect 203250 93550 203252 93602
rect 203196 93044 203252 93550
rect 203196 92978 203252 92988
rect 203980 93042 204036 93660
rect 203980 92990 203982 93042
rect 204034 92990 204036 93042
rect 203980 92978 204036 92990
rect 204316 75572 204372 75582
rect 204316 75478 204372 75516
rect 203980 67060 204036 67070
rect 203196 66946 203252 66958
rect 203196 66894 203198 66946
rect 203250 66894 203252 66946
rect 203196 66836 203252 66894
rect 203196 66770 203252 66780
rect 203980 66386 204036 67004
rect 203980 66334 203982 66386
rect 204034 66334 204036 66386
rect 203980 66322 204036 66334
rect 203756 49922 203812 49934
rect 203756 49870 203758 49922
rect 203810 49870 203812 49922
rect 203756 49364 203812 49870
rect 203756 49298 203812 49308
rect 204092 41298 204148 41310
rect 204092 41246 204094 41298
rect 204146 41246 204148 41298
rect 204092 40628 204148 41246
rect 204092 40562 204148 40572
rect 202412 27682 202468 27692
rect 190652 25330 190708 25340
rect 189456 25116 189720 25126
rect 189512 25060 189560 25116
rect 189616 25060 189664 25116
rect 189456 25050 189720 25060
rect 188796 24332 189060 24342
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 188796 24266 189060 24276
rect 204316 23714 204372 23726
rect 204316 23662 204318 23714
rect 204370 23662 204372 23714
rect 189456 23548 189720 23558
rect 189512 23492 189560 23548
rect 189616 23492 189664 23548
rect 189456 23482 189720 23492
rect 204316 23156 204372 23662
rect 204316 23090 204372 23100
rect 188796 22764 189060 22774
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 188796 22698 189060 22708
rect 189456 21980 189720 21990
rect 189512 21924 189560 21980
rect 189616 21924 189664 21980
rect 189456 21914 189720 21924
rect 188796 21196 189060 21206
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 188796 21130 189060 21140
rect 140028 17054 140030 17106
rect 140082 17054 140084 17106
rect 140028 17042 140084 17054
rect 154364 17108 154420 17118
rect 154588 17108 154644 20412
rect 189456 20412 189720 20422
rect 189512 20356 189560 20412
rect 189616 20356 189664 20412
rect 189456 20346 189720 20356
rect 188796 19628 189060 19638
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 188796 19562 189060 19572
rect 189456 18844 189720 18854
rect 189512 18788 189560 18844
rect 189616 18788 189664 18844
rect 189456 18778 189720 18788
rect 188796 18060 189060 18070
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 188796 17994 189060 18004
rect 158736 17276 159000 17286
rect 158792 17220 158840 17276
rect 158896 17220 158944 17276
rect 158736 17210 159000 17220
rect 189456 17276 189720 17286
rect 189512 17220 189560 17276
rect 189616 17220 189664 17276
rect 189456 17210 189720 17220
rect 154364 17106 154644 17108
rect 154364 17054 154366 17106
rect 154418 17054 154644 17106
rect 154364 17052 154644 17054
rect 154364 17042 154420 17052
rect 67900 16830 67902 16882
rect 67954 16830 67956 16882
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 35856 15708 36120 15718
rect 35912 15652 35960 15708
rect 36016 15652 36064 15708
rect 35856 15642 36120 15652
rect 66576 15708 66840 15718
rect 66632 15652 66680 15708
rect 66736 15652 66784 15708
rect 66576 15642 66840 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 67900 14532 67956 16830
rect 125580 16884 125636 16894
rect 125580 16790 125636 16828
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 127356 16492 127620 16502
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127356 16426 127620 16436
rect 158076 16492 158340 16502
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158076 16426 158340 16436
rect 188796 16492 189060 16502
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 188796 16426 189060 16436
rect 97296 15708 97560 15718
rect 97352 15652 97400 15708
rect 97456 15652 97504 15708
rect 97296 15642 97560 15652
rect 128016 15708 128280 15718
rect 128072 15652 128120 15708
rect 128176 15652 128224 15708
rect 128016 15642 128280 15652
rect 158736 15708 159000 15718
rect 158792 15652 158840 15708
rect 158896 15652 158944 15708
rect 158736 15642 159000 15652
rect 189456 15708 189720 15718
rect 189512 15652 189560 15708
rect 189616 15652 189664 15708
rect 189456 15642 189720 15652
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 127356 14924 127620 14934
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127356 14858 127620 14868
rect 158076 14924 158340 14934
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158076 14858 158340 14868
rect 188796 14924 189060 14934
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 188796 14858 189060 14868
rect 204092 14642 204148 14654
rect 204092 14590 204094 14642
rect 204146 14590 204148 14642
rect 67900 14466 67956 14476
rect 201740 14532 201796 14542
rect 201740 14438 201796 14476
rect 204092 14420 204148 14590
rect 204092 14354 204148 14364
rect 204316 14532 204372 14542
rect 35856 14140 36120 14150
rect 35912 14084 35960 14140
rect 36016 14084 36064 14140
rect 35856 14074 36120 14084
rect 66576 14140 66840 14150
rect 66632 14084 66680 14140
rect 66736 14084 66784 14140
rect 66576 14074 66840 14084
rect 97296 14140 97560 14150
rect 97352 14084 97400 14140
rect 97456 14084 97504 14140
rect 97296 14074 97560 14084
rect 128016 14140 128280 14150
rect 128072 14084 128120 14140
rect 128176 14084 128224 14140
rect 128016 14074 128280 14084
rect 158736 14140 159000 14150
rect 158792 14084 158840 14140
rect 158896 14084 158944 14140
rect 158736 14074 159000 14084
rect 189456 14140 189720 14150
rect 189512 14084 189560 14140
rect 189616 14084 189664 14140
rect 189456 14074 189720 14084
rect 204316 13970 204372 14476
rect 204316 13918 204318 13970
rect 204370 13918 204372 13970
rect 204316 13906 204372 13918
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 127356 13356 127620 13366
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127356 13290 127620 13300
rect 158076 13356 158340 13366
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158076 13290 158340 13300
rect 188796 13356 189060 13366
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 188796 13290 189060 13300
rect 35856 12572 36120 12582
rect 35912 12516 35960 12572
rect 36016 12516 36064 12572
rect 35856 12506 36120 12516
rect 66576 12572 66840 12582
rect 66632 12516 66680 12572
rect 66736 12516 66784 12572
rect 66576 12506 66840 12516
rect 97296 12572 97560 12582
rect 97352 12516 97400 12572
rect 97456 12516 97504 12572
rect 97296 12506 97560 12516
rect 128016 12572 128280 12582
rect 128072 12516 128120 12572
rect 128176 12516 128224 12572
rect 128016 12506 128280 12516
rect 158736 12572 159000 12582
rect 158792 12516 158840 12572
rect 158896 12516 158944 12572
rect 158736 12506 159000 12516
rect 189456 12572 189720 12582
rect 189512 12516 189560 12572
rect 189616 12516 189664 12572
rect 189456 12506 189720 12516
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 127356 11788 127620 11798
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127356 11722 127620 11732
rect 158076 11788 158340 11798
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158076 11722 158340 11732
rect 188796 11788 189060 11798
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 188796 11722 189060 11732
rect 35856 11004 36120 11014
rect 35912 10948 35960 11004
rect 36016 10948 36064 11004
rect 35856 10938 36120 10948
rect 66576 11004 66840 11014
rect 66632 10948 66680 11004
rect 66736 10948 66784 11004
rect 66576 10938 66840 10948
rect 97296 11004 97560 11014
rect 97352 10948 97400 11004
rect 97456 10948 97504 11004
rect 97296 10938 97560 10948
rect 128016 11004 128280 11014
rect 128072 10948 128120 11004
rect 128176 10948 128224 11004
rect 128016 10938 128280 10948
rect 158736 11004 159000 11014
rect 158792 10948 158840 11004
rect 158896 10948 158944 11004
rect 158736 10938 159000 10948
rect 189456 11004 189720 11014
rect 189512 10948 189560 11004
rect 189616 10948 189664 11004
rect 189456 10938 189720 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 127356 10220 127620 10230
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127356 10154 127620 10164
rect 158076 10220 158340 10230
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158076 10154 158340 10164
rect 188796 10220 189060 10230
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 188796 10154 189060 10164
rect 12684 9538 12740 9548
rect 2492 9426 2548 9436
rect 5136 9436 5400 9446
rect 5192 9380 5240 9436
rect 5296 9380 5344 9436
rect 5136 9370 5400 9380
rect 35856 9436 36120 9446
rect 35912 9380 35960 9436
rect 36016 9380 36064 9436
rect 35856 9370 36120 9380
rect 66576 9436 66840 9446
rect 66632 9380 66680 9436
rect 66736 9380 66784 9436
rect 66576 9370 66840 9380
rect 97296 9436 97560 9446
rect 97352 9380 97400 9436
rect 97456 9380 97504 9436
rect 97296 9370 97560 9380
rect 128016 9436 128280 9446
rect 128072 9380 128120 9436
rect 128176 9380 128224 9436
rect 128016 9370 128280 9380
rect 158736 9436 159000 9446
rect 158792 9380 158840 9436
rect 158896 9380 158944 9436
rect 158736 9370 159000 9380
rect 189456 9436 189720 9446
rect 189512 9380 189560 9436
rect 189616 9380 189664 9436
rect 189456 9370 189720 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 127356 8652 127620 8662
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127356 8586 127620 8596
rect 158076 8652 158340 8662
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158076 8586 158340 8596
rect 188796 8652 189060 8662
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 188796 8586 189060 8596
rect 5136 7868 5400 7878
rect 5192 7812 5240 7868
rect 5296 7812 5344 7868
rect 5136 7802 5400 7812
rect 35856 7868 36120 7878
rect 35912 7812 35960 7868
rect 36016 7812 36064 7868
rect 35856 7802 36120 7812
rect 66576 7868 66840 7878
rect 66632 7812 66680 7868
rect 66736 7812 66784 7868
rect 66576 7802 66840 7812
rect 97296 7868 97560 7878
rect 97352 7812 97400 7868
rect 97456 7812 97504 7868
rect 97296 7802 97560 7812
rect 128016 7868 128280 7878
rect 128072 7812 128120 7868
rect 128176 7812 128224 7868
rect 128016 7802 128280 7812
rect 158736 7868 159000 7878
rect 158792 7812 158840 7868
rect 158896 7812 158944 7868
rect 158736 7802 159000 7812
rect 189456 7868 189720 7878
rect 189512 7812 189560 7868
rect 189616 7812 189664 7868
rect 189456 7802 189720 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 127356 7084 127620 7094
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127356 7018 127620 7028
rect 158076 7084 158340 7094
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158076 7018 158340 7028
rect 188796 7084 189060 7094
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 188796 7018 189060 7028
rect 5136 6300 5400 6310
rect 5192 6244 5240 6300
rect 5296 6244 5344 6300
rect 5136 6234 5400 6244
rect 35856 6300 36120 6310
rect 35912 6244 35960 6300
rect 36016 6244 36064 6300
rect 35856 6234 36120 6244
rect 66576 6300 66840 6310
rect 66632 6244 66680 6300
rect 66736 6244 66784 6300
rect 66576 6234 66840 6244
rect 97296 6300 97560 6310
rect 97352 6244 97400 6300
rect 97456 6244 97504 6300
rect 97296 6234 97560 6244
rect 128016 6300 128280 6310
rect 128072 6244 128120 6300
rect 128176 6244 128224 6300
rect 128016 6234 128280 6244
rect 158736 6300 159000 6310
rect 158792 6244 158840 6300
rect 158896 6244 158944 6300
rect 158736 6234 159000 6244
rect 189456 6300 189720 6310
rect 189512 6244 189560 6300
rect 189616 6244 189664 6300
rect 189456 6234 189720 6244
rect 1708 6018 1764 6030
rect 1708 5966 1710 6018
rect 1762 5966 1764 6018
rect 1708 5684 1764 5966
rect 1708 5618 1764 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 127356 5516 127620 5526
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127356 5450 127620 5460
rect 158076 5516 158340 5526
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158076 5450 158340 5460
rect 188796 5516 189060 5526
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 188796 5450 189060 5460
rect 5136 4732 5400 4742
rect 5192 4676 5240 4732
rect 5296 4676 5344 4732
rect 5136 4666 5400 4676
rect 35856 4732 36120 4742
rect 35912 4676 35960 4732
rect 36016 4676 36064 4732
rect 35856 4666 36120 4676
rect 66576 4732 66840 4742
rect 66632 4676 66680 4732
rect 66736 4676 66784 4732
rect 66576 4666 66840 4676
rect 97296 4732 97560 4742
rect 97352 4676 97400 4732
rect 97456 4676 97504 4732
rect 97296 4666 97560 4676
rect 128016 4732 128280 4742
rect 128072 4676 128120 4732
rect 128176 4676 128224 4732
rect 128016 4666 128280 4676
rect 158736 4732 159000 4742
rect 158792 4676 158840 4732
rect 158896 4676 158944 4732
rect 158736 4666 159000 4676
rect 189456 4732 189720 4742
rect 189512 4676 189560 4732
rect 189616 4676 189664 4732
rect 189456 4666 189720 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 127356 3948 127620 3958
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127356 3882 127620 3892
rect 158076 3948 158340 3958
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158076 3882 158340 3892
rect 188796 3948 189060 3958
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 188796 3882 189060 3892
rect 1708 3666 1764 3678
rect 1708 3614 1710 3666
rect 1762 3614 1764 3666
rect 1708 1876 1764 3614
rect 34524 3332 34580 3342
rect 103068 3332 103124 3342
rect 171612 3332 171668 3342
rect 34300 3330 34580 3332
rect 34300 3278 34526 3330
rect 34578 3278 34580 3330
rect 34300 3276 34580 3278
rect 5136 3164 5400 3174
rect 5192 3108 5240 3164
rect 5296 3108 5344 3164
rect 5136 3098 5400 3108
rect 1708 1810 1764 1820
rect 34300 800 34356 3276
rect 34524 3266 34580 3276
rect 102844 3330 103124 3332
rect 102844 3278 103070 3330
rect 103122 3278 103124 3330
rect 102844 3276 103124 3278
rect 35856 3164 36120 3174
rect 35912 3108 35960 3164
rect 36016 3108 36064 3164
rect 35856 3098 36120 3108
rect 66576 3164 66840 3174
rect 66632 3108 66680 3164
rect 66736 3108 66784 3164
rect 66576 3098 66840 3108
rect 97296 3164 97560 3174
rect 97352 3108 97400 3164
rect 97456 3108 97504 3164
rect 97296 3098 97560 3108
rect 102844 800 102900 3276
rect 103068 3266 103124 3276
rect 171388 3330 171668 3332
rect 171388 3278 171614 3330
rect 171666 3278 171668 3330
rect 171388 3276 171668 3278
rect 128016 3164 128280 3174
rect 128072 3108 128120 3164
rect 128176 3108 128224 3164
rect 128016 3098 128280 3108
rect 158736 3164 159000 3174
rect 158792 3108 158840 3164
rect 158896 3108 158944 3164
rect 158736 3098 159000 3108
rect 171388 800 171444 3276
rect 171612 3266 171668 3276
rect 189456 3164 189720 3174
rect 189512 3108 189560 3164
rect 189616 3108 189664 3164
rect 189456 3098 189720 3108
rect 34272 0 34384 800
rect 102816 0 102928 800
rect 171360 0 171472 800
<< via2 >>
rect 1708 157836 1764 157892
rect 1708 154140 1764 154196
rect 1708 150332 1764 150388
rect 1820 146524 1876 146580
rect 1708 142716 1764 142772
rect 1708 138962 1764 138964
rect 1708 138910 1710 138962
rect 1710 138910 1762 138962
rect 1762 138910 1764 138962
rect 1708 138908 1764 138910
rect 1708 135100 1764 135156
rect 1708 131292 1764 131348
rect 1708 127484 1764 127540
rect 1820 123730 1876 123732
rect 1820 123678 1822 123730
rect 1822 123678 1874 123730
rect 1874 123678 1876 123730
rect 1820 123676 1876 123678
rect 1708 119868 1764 119924
rect 1708 116060 1764 116116
rect 1708 112252 1764 112308
rect 1708 108498 1764 108500
rect 1708 108446 1710 108498
rect 1710 108446 1762 108498
rect 1762 108446 1764 108498
rect 1708 108444 1764 108446
rect 1708 104636 1764 104692
rect 2044 101666 2100 101668
rect 2044 101614 2046 101666
rect 2046 101614 2098 101666
rect 2098 101614 2100 101666
rect 2044 101612 2100 101614
rect 1708 101388 1764 101444
rect 1708 100828 1764 100884
rect 1708 97020 1764 97076
rect 1708 93490 1764 93492
rect 1708 93438 1710 93490
rect 1710 93438 1762 93490
rect 1762 93438 1764 93490
rect 1708 93436 1764 93438
rect 1708 89404 1764 89460
rect 1708 85596 1764 85652
rect 1708 82066 1764 82068
rect 1708 82014 1710 82066
rect 1710 82014 1762 82066
rect 1762 82014 1764 82066
rect 1708 82012 1764 82014
rect 1708 78594 1764 78596
rect 1708 78542 1710 78594
rect 1710 78542 1762 78594
rect 1762 78542 1764 78594
rect 1708 78540 1764 78542
rect 1708 77980 1764 78036
rect 2044 75628 2100 75684
rect 2156 74732 2212 74788
rect 2268 76300 2324 76356
rect 1708 74172 1764 74228
rect 1708 70364 1764 70420
rect 1708 66556 1764 66612
rect 1708 62914 1764 62916
rect 1708 62862 1710 62914
rect 1710 62862 1762 62914
rect 1762 62862 1764 62914
rect 1708 62860 1764 62862
rect 1708 58994 1764 58996
rect 1708 58942 1710 58994
rect 1710 58942 1762 58994
rect 1762 58942 1764 58994
rect 1708 58940 1764 58942
rect 2268 55298 2324 55300
rect 2268 55246 2270 55298
rect 2270 55246 2322 55298
rect 2322 55246 2324 55298
rect 2268 55244 2324 55246
rect 1708 55186 1764 55188
rect 1708 55134 1710 55186
rect 1710 55134 1762 55186
rect 1762 55134 1764 55186
rect 1708 55132 1764 55134
rect 1708 51324 1764 51380
rect 1708 47516 1764 47572
rect 2268 44322 2324 44324
rect 2268 44270 2270 44322
rect 2270 44270 2322 44322
rect 2322 44270 2324 44322
rect 2268 44268 2324 44270
rect 1820 43762 1876 43764
rect 1820 43710 1822 43762
rect 1822 43710 1874 43762
rect 1874 43710 1876 43762
rect 1820 43708 1876 43710
rect 1708 39900 1764 39956
rect 1708 36092 1764 36148
rect 2044 36204 2100 36260
rect 2156 34636 2212 34692
rect 1708 32284 1764 32340
rect 1708 28530 1764 28532
rect 1708 28478 1710 28530
rect 1710 28478 1762 28530
rect 1762 28478 1764 28530
rect 1708 28476 1764 28478
rect 1708 24668 1764 24724
rect 5136 156826 5192 156828
rect 5136 156774 5138 156826
rect 5138 156774 5190 156826
rect 5190 156774 5192 156826
rect 5136 156772 5192 156774
rect 5240 156826 5296 156828
rect 5240 156774 5242 156826
rect 5242 156774 5294 156826
rect 5294 156774 5296 156826
rect 5240 156772 5296 156774
rect 5344 156826 5400 156828
rect 5344 156774 5346 156826
rect 5346 156774 5398 156826
rect 5398 156774 5400 156826
rect 5344 156772 5400 156774
rect 20076 156322 20132 156324
rect 20076 156270 20078 156322
rect 20078 156270 20130 156322
rect 20130 156270 20132 156322
rect 20076 156268 20132 156270
rect 22764 156268 22820 156324
rect 4476 156042 4532 156044
rect 4476 155990 4478 156042
rect 4478 155990 4530 156042
rect 4530 155990 4532 156042
rect 4476 155988 4532 155990
rect 4580 156042 4636 156044
rect 4580 155990 4582 156042
rect 4582 155990 4634 156042
rect 4634 155990 4636 156042
rect 4580 155988 4636 155990
rect 4684 156042 4740 156044
rect 4684 155990 4686 156042
rect 4686 155990 4738 156042
rect 4738 155990 4740 156042
rect 4684 155988 4740 155990
rect 5136 155258 5192 155260
rect 5136 155206 5138 155258
rect 5138 155206 5190 155258
rect 5190 155206 5192 155258
rect 5136 155204 5192 155206
rect 5240 155258 5296 155260
rect 5240 155206 5242 155258
rect 5242 155206 5294 155258
rect 5294 155206 5296 155258
rect 5240 155204 5296 155206
rect 5344 155258 5400 155260
rect 5344 155206 5346 155258
rect 5346 155206 5398 155258
rect 5398 155206 5400 155258
rect 5344 155204 5400 155206
rect 4476 154474 4532 154476
rect 4476 154422 4478 154474
rect 4478 154422 4530 154474
rect 4530 154422 4532 154474
rect 4476 154420 4532 154422
rect 4580 154474 4636 154476
rect 4580 154422 4582 154474
rect 4582 154422 4634 154474
rect 4634 154422 4636 154474
rect 4580 154420 4636 154422
rect 4684 154474 4740 154476
rect 4684 154422 4686 154474
rect 4686 154422 4738 154474
rect 4738 154422 4740 154474
rect 4684 154420 4740 154422
rect 5136 153690 5192 153692
rect 5136 153638 5138 153690
rect 5138 153638 5190 153690
rect 5190 153638 5192 153690
rect 5136 153636 5192 153638
rect 5240 153690 5296 153692
rect 5240 153638 5242 153690
rect 5242 153638 5294 153690
rect 5294 153638 5296 153690
rect 5240 153636 5296 153638
rect 5344 153690 5400 153692
rect 5344 153638 5346 153690
rect 5346 153638 5398 153690
rect 5398 153638 5400 153690
rect 5344 153636 5400 153638
rect 4476 152906 4532 152908
rect 4476 152854 4478 152906
rect 4478 152854 4530 152906
rect 4530 152854 4532 152906
rect 4476 152852 4532 152854
rect 4580 152906 4636 152908
rect 4580 152854 4582 152906
rect 4582 152854 4634 152906
rect 4634 152854 4636 152906
rect 4580 152852 4636 152854
rect 4684 152906 4740 152908
rect 4684 152854 4686 152906
rect 4686 152854 4738 152906
rect 4738 152854 4740 152906
rect 4684 152852 4740 152854
rect 5136 152122 5192 152124
rect 5136 152070 5138 152122
rect 5138 152070 5190 152122
rect 5190 152070 5192 152122
rect 5136 152068 5192 152070
rect 5240 152122 5296 152124
rect 5240 152070 5242 152122
rect 5242 152070 5294 152122
rect 5294 152070 5296 152122
rect 5240 152068 5296 152070
rect 5344 152122 5400 152124
rect 5344 152070 5346 152122
rect 5346 152070 5398 152122
rect 5398 152070 5400 152122
rect 5344 152068 5400 152070
rect 4476 151338 4532 151340
rect 4476 151286 4478 151338
rect 4478 151286 4530 151338
rect 4530 151286 4532 151338
rect 4476 151284 4532 151286
rect 4580 151338 4636 151340
rect 4580 151286 4582 151338
rect 4582 151286 4634 151338
rect 4634 151286 4636 151338
rect 4580 151284 4636 151286
rect 4684 151338 4740 151340
rect 4684 151286 4686 151338
rect 4686 151286 4738 151338
rect 4738 151286 4740 151338
rect 4684 151284 4740 151286
rect 5136 150554 5192 150556
rect 5136 150502 5138 150554
rect 5138 150502 5190 150554
rect 5190 150502 5192 150554
rect 5136 150500 5192 150502
rect 5240 150554 5296 150556
rect 5240 150502 5242 150554
rect 5242 150502 5294 150554
rect 5294 150502 5296 150554
rect 5240 150500 5296 150502
rect 5344 150554 5400 150556
rect 5344 150502 5346 150554
rect 5346 150502 5398 150554
rect 5398 150502 5400 150554
rect 5344 150500 5400 150502
rect 4476 149770 4532 149772
rect 4476 149718 4478 149770
rect 4478 149718 4530 149770
rect 4530 149718 4532 149770
rect 4476 149716 4532 149718
rect 4580 149770 4636 149772
rect 4580 149718 4582 149770
rect 4582 149718 4634 149770
rect 4634 149718 4636 149770
rect 4580 149716 4636 149718
rect 4684 149770 4740 149772
rect 4684 149718 4686 149770
rect 4686 149718 4738 149770
rect 4738 149718 4740 149770
rect 4684 149716 4740 149718
rect 5136 148986 5192 148988
rect 5136 148934 5138 148986
rect 5138 148934 5190 148986
rect 5190 148934 5192 148986
rect 5136 148932 5192 148934
rect 5240 148986 5296 148988
rect 5240 148934 5242 148986
rect 5242 148934 5294 148986
rect 5294 148934 5296 148986
rect 5240 148932 5296 148934
rect 5344 148986 5400 148988
rect 5344 148934 5346 148986
rect 5346 148934 5398 148986
rect 5398 148934 5400 148986
rect 5344 148932 5400 148934
rect 4476 148202 4532 148204
rect 4476 148150 4478 148202
rect 4478 148150 4530 148202
rect 4530 148150 4532 148202
rect 4476 148148 4532 148150
rect 4580 148202 4636 148204
rect 4580 148150 4582 148202
rect 4582 148150 4634 148202
rect 4634 148150 4636 148202
rect 4580 148148 4636 148150
rect 4684 148202 4740 148204
rect 4684 148150 4686 148202
rect 4686 148150 4738 148202
rect 4738 148150 4740 148202
rect 4684 148148 4740 148150
rect 5136 147418 5192 147420
rect 5136 147366 5138 147418
rect 5138 147366 5190 147418
rect 5190 147366 5192 147418
rect 5136 147364 5192 147366
rect 5240 147418 5296 147420
rect 5240 147366 5242 147418
rect 5242 147366 5294 147418
rect 5294 147366 5296 147418
rect 5240 147364 5296 147366
rect 5344 147418 5400 147420
rect 5344 147366 5346 147418
rect 5346 147366 5398 147418
rect 5398 147366 5400 147418
rect 5344 147364 5400 147366
rect 2828 146914 2884 146916
rect 2828 146862 2830 146914
rect 2830 146862 2882 146914
rect 2882 146862 2884 146914
rect 2828 146860 2884 146862
rect 12572 146860 12628 146916
rect 4476 146634 4532 146636
rect 4476 146582 4478 146634
rect 4478 146582 4530 146634
rect 4530 146582 4532 146634
rect 4476 146580 4532 146582
rect 4580 146634 4636 146636
rect 4580 146582 4582 146634
rect 4582 146582 4634 146634
rect 4634 146582 4636 146634
rect 4580 146580 4636 146582
rect 4684 146634 4740 146636
rect 4684 146582 4686 146634
rect 4686 146582 4738 146634
rect 4738 146582 4740 146634
rect 4684 146580 4740 146582
rect 5136 145850 5192 145852
rect 5136 145798 5138 145850
rect 5138 145798 5190 145850
rect 5190 145798 5192 145850
rect 5136 145796 5192 145798
rect 5240 145850 5296 145852
rect 5240 145798 5242 145850
rect 5242 145798 5294 145850
rect 5294 145798 5296 145850
rect 5240 145796 5296 145798
rect 5344 145850 5400 145852
rect 5344 145798 5346 145850
rect 5346 145798 5398 145850
rect 5398 145798 5400 145850
rect 5344 145796 5400 145798
rect 4476 145066 4532 145068
rect 4476 145014 4478 145066
rect 4478 145014 4530 145066
rect 4530 145014 4532 145066
rect 4476 145012 4532 145014
rect 4580 145066 4636 145068
rect 4580 145014 4582 145066
rect 4582 145014 4634 145066
rect 4634 145014 4636 145066
rect 4580 145012 4636 145014
rect 4684 145066 4740 145068
rect 4684 145014 4686 145066
rect 4686 145014 4738 145066
rect 4738 145014 4740 145066
rect 4684 145012 4740 145014
rect 5136 144282 5192 144284
rect 5136 144230 5138 144282
rect 5138 144230 5190 144282
rect 5190 144230 5192 144282
rect 5136 144228 5192 144230
rect 5240 144282 5296 144284
rect 5240 144230 5242 144282
rect 5242 144230 5294 144282
rect 5294 144230 5296 144282
rect 5240 144228 5296 144230
rect 5344 144282 5400 144284
rect 5344 144230 5346 144282
rect 5346 144230 5398 144282
rect 5398 144230 5400 144282
rect 5344 144228 5400 144230
rect 4476 143498 4532 143500
rect 4476 143446 4478 143498
rect 4478 143446 4530 143498
rect 4530 143446 4532 143498
rect 4476 143444 4532 143446
rect 4580 143498 4636 143500
rect 4580 143446 4582 143498
rect 4582 143446 4634 143498
rect 4634 143446 4636 143498
rect 4580 143444 4636 143446
rect 4684 143498 4740 143500
rect 4684 143446 4686 143498
rect 4686 143446 4738 143498
rect 4738 143446 4740 143498
rect 4684 143444 4740 143446
rect 5136 142714 5192 142716
rect 5136 142662 5138 142714
rect 5138 142662 5190 142714
rect 5190 142662 5192 142714
rect 5136 142660 5192 142662
rect 5240 142714 5296 142716
rect 5240 142662 5242 142714
rect 5242 142662 5294 142714
rect 5294 142662 5296 142714
rect 5240 142660 5296 142662
rect 5344 142714 5400 142716
rect 5344 142662 5346 142714
rect 5346 142662 5398 142714
rect 5398 142662 5400 142714
rect 5344 142660 5400 142662
rect 4476 141930 4532 141932
rect 4476 141878 4478 141930
rect 4478 141878 4530 141930
rect 4530 141878 4532 141930
rect 4476 141876 4532 141878
rect 4580 141930 4636 141932
rect 4580 141878 4582 141930
rect 4582 141878 4634 141930
rect 4634 141878 4636 141930
rect 4580 141876 4636 141878
rect 4684 141930 4740 141932
rect 4684 141878 4686 141930
rect 4686 141878 4738 141930
rect 4738 141878 4740 141930
rect 4684 141876 4740 141878
rect 5136 141146 5192 141148
rect 5136 141094 5138 141146
rect 5138 141094 5190 141146
rect 5190 141094 5192 141146
rect 5136 141092 5192 141094
rect 5240 141146 5296 141148
rect 5240 141094 5242 141146
rect 5242 141094 5294 141146
rect 5294 141094 5296 141146
rect 5240 141092 5296 141094
rect 5344 141146 5400 141148
rect 5344 141094 5346 141146
rect 5346 141094 5398 141146
rect 5398 141094 5400 141146
rect 5344 141092 5400 141094
rect 4476 140362 4532 140364
rect 4476 140310 4478 140362
rect 4478 140310 4530 140362
rect 4530 140310 4532 140362
rect 4476 140308 4532 140310
rect 4580 140362 4636 140364
rect 4580 140310 4582 140362
rect 4582 140310 4634 140362
rect 4634 140310 4636 140362
rect 4580 140308 4636 140310
rect 4684 140362 4740 140364
rect 4684 140310 4686 140362
rect 4686 140310 4738 140362
rect 4738 140310 4740 140362
rect 4684 140308 4740 140310
rect 5136 139578 5192 139580
rect 5136 139526 5138 139578
rect 5138 139526 5190 139578
rect 5190 139526 5192 139578
rect 5136 139524 5192 139526
rect 5240 139578 5296 139580
rect 5240 139526 5242 139578
rect 5242 139526 5294 139578
rect 5294 139526 5296 139578
rect 5240 139524 5296 139526
rect 5344 139578 5400 139580
rect 5344 139526 5346 139578
rect 5346 139526 5398 139578
rect 5398 139526 5400 139578
rect 5344 139524 5400 139526
rect 4476 138794 4532 138796
rect 4476 138742 4478 138794
rect 4478 138742 4530 138794
rect 4530 138742 4532 138794
rect 4476 138740 4532 138742
rect 4580 138794 4636 138796
rect 4580 138742 4582 138794
rect 4582 138742 4634 138794
rect 4634 138742 4636 138794
rect 4580 138740 4636 138742
rect 4684 138794 4740 138796
rect 4684 138742 4686 138794
rect 4686 138742 4738 138794
rect 4738 138742 4740 138794
rect 4684 138740 4740 138742
rect 5136 138010 5192 138012
rect 5136 137958 5138 138010
rect 5138 137958 5190 138010
rect 5190 137958 5192 138010
rect 5136 137956 5192 137958
rect 5240 138010 5296 138012
rect 5240 137958 5242 138010
rect 5242 137958 5294 138010
rect 5294 137958 5296 138010
rect 5240 137956 5296 137958
rect 5344 138010 5400 138012
rect 5344 137958 5346 138010
rect 5346 137958 5398 138010
rect 5398 137958 5400 138010
rect 5344 137956 5400 137958
rect 4476 137226 4532 137228
rect 4476 137174 4478 137226
rect 4478 137174 4530 137226
rect 4530 137174 4532 137226
rect 4476 137172 4532 137174
rect 4580 137226 4636 137228
rect 4580 137174 4582 137226
rect 4582 137174 4634 137226
rect 4634 137174 4636 137226
rect 4580 137172 4636 137174
rect 4684 137226 4740 137228
rect 4684 137174 4686 137226
rect 4686 137174 4738 137226
rect 4738 137174 4740 137226
rect 4684 137172 4740 137174
rect 5136 136442 5192 136444
rect 5136 136390 5138 136442
rect 5138 136390 5190 136442
rect 5190 136390 5192 136442
rect 5136 136388 5192 136390
rect 5240 136442 5296 136444
rect 5240 136390 5242 136442
rect 5242 136390 5294 136442
rect 5294 136390 5296 136442
rect 5240 136388 5296 136390
rect 5344 136442 5400 136444
rect 5344 136390 5346 136442
rect 5346 136390 5398 136442
rect 5398 136390 5400 136442
rect 5344 136388 5400 136390
rect 4476 135658 4532 135660
rect 4476 135606 4478 135658
rect 4478 135606 4530 135658
rect 4530 135606 4532 135658
rect 4476 135604 4532 135606
rect 4580 135658 4636 135660
rect 4580 135606 4582 135658
rect 4582 135606 4634 135658
rect 4634 135606 4636 135658
rect 4580 135604 4636 135606
rect 4684 135658 4740 135660
rect 4684 135606 4686 135658
rect 4686 135606 4738 135658
rect 4738 135606 4740 135658
rect 4684 135604 4740 135606
rect 2828 135154 2884 135156
rect 2828 135102 2830 135154
rect 2830 135102 2882 135154
rect 2882 135102 2884 135154
rect 2828 135100 2884 135102
rect 5136 134874 5192 134876
rect 5136 134822 5138 134874
rect 5138 134822 5190 134874
rect 5190 134822 5192 134874
rect 5136 134820 5192 134822
rect 5240 134874 5296 134876
rect 5240 134822 5242 134874
rect 5242 134822 5294 134874
rect 5294 134822 5296 134874
rect 5240 134820 5296 134822
rect 5344 134874 5400 134876
rect 5344 134822 5346 134874
rect 5346 134822 5398 134874
rect 5398 134822 5400 134874
rect 5344 134820 5400 134822
rect 4476 134090 4532 134092
rect 4476 134038 4478 134090
rect 4478 134038 4530 134090
rect 4530 134038 4532 134090
rect 4476 134036 4532 134038
rect 4580 134090 4636 134092
rect 4580 134038 4582 134090
rect 4582 134038 4634 134090
rect 4634 134038 4636 134090
rect 4580 134036 4636 134038
rect 4684 134090 4740 134092
rect 4684 134038 4686 134090
rect 4686 134038 4738 134090
rect 4738 134038 4740 134090
rect 4684 134036 4740 134038
rect 5136 133306 5192 133308
rect 5136 133254 5138 133306
rect 5138 133254 5190 133306
rect 5190 133254 5192 133306
rect 5136 133252 5192 133254
rect 5240 133306 5296 133308
rect 5240 133254 5242 133306
rect 5242 133254 5294 133306
rect 5294 133254 5296 133306
rect 5240 133252 5296 133254
rect 5344 133306 5400 133308
rect 5344 133254 5346 133306
rect 5346 133254 5398 133306
rect 5398 133254 5400 133306
rect 5344 133252 5400 133254
rect 4476 132522 4532 132524
rect 4476 132470 4478 132522
rect 4478 132470 4530 132522
rect 4530 132470 4532 132522
rect 4476 132468 4532 132470
rect 4580 132522 4636 132524
rect 4580 132470 4582 132522
rect 4582 132470 4634 132522
rect 4634 132470 4636 132522
rect 4580 132468 4636 132470
rect 4684 132522 4740 132524
rect 4684 132470 4686 132522
rect 4686 132470 4738 132522
rect 4738 132470 4740 132522
rect 4684 132468 4740 132470
rect 5136 131738 5192 131740
rect 5136 131686 5138 131738
rect 5138 131686 5190 131738
rect 5190 131686 5192 131738
rect 5136 131684 5192 131686
rect 5240 131738 5296 131740
rect 5240 131686 5242 131738
rect 5242 131686 5294 131738
rect 5294 131686 5296 131738
rect 5240 131684 5296 131686
rect 5344 131738 5400 131740
rect 5344 131686 5346 131738
rect 5346 131686 5398 131738
rect 5398 131686 5400 131738
rect 5344 131684 5400 131686
rect 4476 130954 4532 130956
rect 4476 130902 4478 130954
rect 4478 130902 4530 130954
rect 4530 130902 4532 130954
rect 4476 130900 4532 130902
rect 4580 130954 4636 130956
rect 4580 130902 4582 130954
rect 4582 130902 4634 130954
rect 4634 130902 4636 130954
rect 4580 130900 4636 130902
rect 4684 130954 4740 130956
rect 4684 130902 4686 130954
rect 4686 130902 4738 130954
rect 4738 130902 4740 130954
rect 4684 130900 4740 130902
rect 5136 130170 5192 130172
rect 5136 130118 5138 130170
rect 5138 130118 5190 130170
rect 5190 130118 5192 130170
rect 5136 130116 5192 130118
rect 5240 130170 5296 130172
rect 5240 130118 5242 130170
rect 5242 130118 5294 130170
rect 5294 130118 5296 130170
rect 5240 130116 5296 130118
rect 5344 130170 5400 130172
rect 5344 130118 5346 130170
rect 5346 130118 5398 130170
rect 5398 130118 5400 130170
rect 5344 130116 5400 130118
rect 4476 129386 4532 129388
rect 4476 129334 4478 129386
rect 4478 129334 4530 129386
rect 4530 129334 4532 129386
rect 4476 129332 4532 129334
rect 4580 129386 4636 129388
rect 4580 129334 4582 129386
rect 4582 129334 4634 129386
rect 4634 129334 4636 129386
rect 4580 129332 4636 129334
rect 4684 129386 4740 129388
rect 4684 129334 4686 129386
rect 4686 129334 4738 129386
rect 4738 129334 4740 129386
rect 4684 129332 4740 129334
rect 5136 128602 5192 128604
rect 5136 128550 5138 128602
rect 5138 128550 5190 128602
rect 5190 128550 5192 128602
rect 5136 128548 5192 128550
rect 5240 128602 5296 128604
rect 5240 128550 5242 128602
rect 5242 128550 5294 128602
rect 5294 128550 5296 128602
rect 5240 128548 5296 128550
rect 5344 128602 5400 128604
rect 5344 128550 5346 128602
rect 5346 128550 5398 128602
rect 5398 128550 5400 128602
rect 5344 128548 5400 128550
rect 4476 127818 4532 127820
rect 4476 127766 4478 127818
rect 4478 127766 4530 127818
rect 4530 127766 4532 127818
rect 4476 127764 4532 127766
rect 4580 127818 4636 127820
rect 4580 127766 4582 127818
rect 4582 127766 4634 127818
rect 4634 127766 4636 127818
rect 4580 127764 4636 127766
rect 4684 127818 4740 127820
rect 4684 127766 4686 127818
rect 4686 127766 4738 127818
rect 4738 127766 4740 127818
rect 4684 127764 4740 127766
rect 5136 127034 5192 127036
rect 5136 126982 5138 127034
rect 5138 126982 5190 127034
rect 5190 126982 5192 127034
rect 5136 126980 5192 126982
rect 5240 127034 5296 127036
rect 5240 126982 5242 127034
rect 5242 126982 5294 127034
rect 5294 126982 5296 127034
rect 5240 126980 5296 126982
rect 5344 127034 5400 127036
rect 5344 126982 5346 127034
rect 5346 126982 5398 127034
rect 5398 126982 5400 127034
rect 5344 126980 5400 126982
rect 4476 126250 4532 126252
rect 4476 126198 4478 126250
rect 4478 126198 4530 126250
rect 4530 126198 4532 126250
rect 4476 126196 4532 126198
rect 4580 126250 4636 126252
rect 4580 126198 4582 126250
rect 4582 126198 4634 126250
rect 4634 126198 4636 126250
rect 4580 126196 4636 126198
rect 4684 126250 4740 126252
rect 4684 126198 4686 126250
rect 4686 126198 4738 126250
rect 4738 126198 4740 126250
rect 4684 126196 4740 126198
rect 5136 125466 5192 125468
rect 5136 125414 5138 125466
rect 5138 125414 5190 125466
rect 5190 125414 5192 125466
rect 5136 125412 5192 125414
rect 5240 125466 5296 125468
rect 5240 125414 5242 125466
rect 5242 125414 5294 125466
rect 5294 125414 5296 125466
rect 5240 125412 5296 125414
rect 5344 125466 5400 125468
rect 5344 125414 5346 125466
rect 5346 125414 5398 125466
rect 5398 125414 5400 125466
rect 5344 125412 5400 125414
rect 4476 124682 4532 124684
rect 4476 124630 4478 124682
rect 4478 124630 4530 124682
rect 4530 124630 4532 124682
rect 4476 124628 4532 124630
rect 4580 124682 4636 124684
rect 4580 124630 4582 124682
rect 4582 124630 4634 124682
rect 4634 124630 4636 124682
rect 4580 124628 4636 124630
rect 4684 124682 4740 124684
rect 4684 124630 4686 124682
rect 4686 124630 4738 124682
rect 4738 124630 4740 124682
rect 4684 124628 4740 124630
rect 2828 124178 2884 124180
rect 2828 124126 2830 124178
rect 2830 124126 2882 124178
rect 2882 124126 2884 124178
rect 2828 124124 2884 124126
rect 5136 123898 5192 123900
rect 5136 123846 5138 123898
rect 5138 123846 5190 123898
rect 5190 123846 5192 123898
rect 5136 123844 5192 123846
rect 5240 123898 5296 123900
rect 5240 123846 5242 123898
rect 5242 123846 5294 123898
rect 5294 123846 5296 123898
rect 5240 123844 5296 123846
rect 5344 123898 5400 123900
rect 5344 123846 5346 123898
rect 5346 123846 5398 123898
rect 5398 123846 5400 123898
rect 5344 123844 5400 123846
rect 4476 123114 4532 123116
rect 4476 123062 4478 123114
rect 4478 123062 4530 123114
rect 4530 123062 4532 123114
rect 4476 123060 4532 123062
rect 4580 123114 4636 123116
rect 4580 123062 4582 123114
rect 4582 123062 4634 123114
rect 4634 123062 4636 123114
rect 4580 123060 4636 123062
rect 4684 123114 4740 123116
rect 4684 123062 4686 123114
rect 4686 123062 4738 123114
rect 4738 123062 4740 123114
rect 4684 123060 4740 123062
rect 5136 122330 5192 122332
rect 5136 122278 5138 122330
rect 5138 122278 5190 122330
rect 5190 122278 5192 122330
rect 5136 122276 5192 122278
rect 5240 122330 5296 122332
rect 5240 122278 5242 122330
rect 5242 122278 5294 122330
rect 5294 122278 5296 122330
rect 5240 122276 5296 122278
rect 5344 122330 5400 122332
rect 5344 122278 5346 122330
rect 5346 122278 5398 122330
rect 5398 122278 5400 122330
rect 5344 122276 5400 122278
rect 4476 121546 4532 121548
rect 4476 121494 4478 121546
rect 4478 121494 4530 121546
rect 4530 121494 4532 121546
rect 4476 121492 4532 121494
rect 4580 121546 4636 121548
rect 4580 121494 4582 121546
rect 4582 121494 4634 121546
rect 4634 121494 4636 121546
rect 4580 121492 4636 121494
rect 4684 121546 4740 121548
rect 4684 121494 4686 121546
rect 4686 121494 4738 121546
rect 4738 121494 4740 121546
rect 4684 121492 4740 121494
rect 5136 120762 5192 120764
rect 5136 120710 5138 120762
rect 5138 120710 5190 120762
rect 5190 120710 5192 120762
rect 5136 120708 5192 120710
rect 5240 120762 5296 120764
rect 5240 120710 5242 120762
rect 5242 120710 5294 120762
rect 5294 120710 5296 120762
rect 5240 120708 5296 120710
rect 5344 120762 5400 120764
rect 5344 120710 5346 120762
rect 5346 120710 5398 120762
rect 5398 120710 5400 120762
rect 5344 120708 5400 120710
rect 4476 119978 4532 119980
rect 4476 119926 4478 119978
rect 4478 119926 4530 119978
rect 4530 119926 4532 119978
rect 4476 119924 4532 119926
rect 4580 119978 4636 119980
rect 4580 119926 4582 119978
rect 4582 119926 4634 119978
rect 4634 119926 4636 119978
rect 4580 119924 4636 119926
rect 4684 119978 4740 119980
rect 4684 119926 4686 119978
rect 4686 119926 4738 119978
rect 4738 119926 4740 119978
rect 4684 119924 4740 119926
rect 5136 119194 5192 119196
rect 5136 119142 5138 119194
rect 5138 119142 5190 119194
rect 5190 119142 5192 119194
rect 5136 119140 5192 119142
rect 5240 119194 5296 119196
rect 5240 119142 5242 119194
rect 5242 119142 5294 119194
rect 5294 119142 5296 119194
rect 5240 119140 5296 119142
rect 5344 119194 5400 119196
rect 5344 119142 5346 119194
rect 5346 119142 5398 119194
rect 5398 119142 5400 119194
rect 5344 119140 5400 119142
rect 4476 118410 4532 118412
rect 4476 118358 4478 118410
rect 4478 118358 4530 118410
rect 4530 118358 4532 118410
rect 4476 118356 4532 118358
rect 4580 118410 4636 118412
rect 4580 118358 4582 118410
rect 4582 118358 4634 118410
rect 4634 118358 4636 118410
rect 4580 118356 4636 118358
rect 4684 118410 4740 118412
rect 4684 118358 4686 118410
rect 4686 118358 4738 118410
rect 4738 118358 4740 118410
rect 4684 118356 4740 118358
rect 5136 117626 5192 117628
rect 5136 117574 5138 117626
rect 5138 117574 5190 117626
rect 5190 117574 5192 117626
rect 5136 117572 5192 117574
rect 5240 117626 5296 117628
rect 5240 117574 5242 117626
rect 5242 117574 5294 117626
rect 5294 117574 5296 117626
rect 5240 117572 5296 117574
rect 5344 117626 5400 117628
rect 5344 117574 5346 117626
rect 5346 117574 5398 117626
rect 5398 117574 5400 117626
rect 5344 117572 5400 117574
rect 4476 116842 4532 116844
rect 4476 116790 4478 116842
rect 4478 116790 4530 116842
rect 4530 116790 4532 116842
rect 4476 116788 4532 116790
rect 4580 116842 4636 116844
rect 4580 116790 4582 116842
rect 4582 116790 4634 116842
rect 4634 116790 4636 116842
rect 4580 116788 4636 116790
rect 4684 116842 4740 116844
rect 4684 116790 4686 116842
rect 4686 116790 4738 116842
rect 4738 116790 4740 116842
rect 4684 116788 4740 116790
rect 5136 116058 5192 116060
rect 5136 116006 5138 116058
rect 5138 116006 5190 116058
rect 5190 116006 5192 116058
rect 5136 116004 5192 116006
rect 5240 116058 5296 116060
rect 5240 116006 5242 116058
rect 5242 116006 5294 116058
rect 5294 116006 5296 116058
rect 5240 116004 5296 116006
rect 5344 116058 5400 116060
rect 5344 116006 5346 116058
rect 5346 116006 5398 116058
rect 5398 116006 5400 116058
rect 5344 116004 5400 116006
rect 4476 115274 4532 115276
rect 4476 115222 4478 115274
rect 4478 115222 4530 115274
rect 4530 115222 4532 115274
rect 4476 115220 4532 115222
rect 4580 115274 4636 115276
rect 4580 115222 4582 115274
rect 4582 115222 4634 115274
rect 4634 115222 4636 115274
rect 4580 115220 4636 115222
rect 4684 115274 4740 115276
rect 4684 115222 4686 115274
rect 4686 115222 4738 115274
rect 4738 115222 4740 115274
rect 4684 115220 4740 115222
rect 5136 114490 5192 114492
rect 5136 114438 5138 114490
rect 5138 114438 5190 114490
rect 5190 114438 5192 114490
rect 5136 114436 5192 114438
rect 5240 114490 5296 114492
rect 5240 114438 5242 114490
rect 5242 114438 5294 114490
rect 5294 114438 5296 114490
rect 5240 114436 5296 114438
rect 5344 114490 5400 114492
rect 5344 114438 5346 114490
rect 5346 114438 5398 114490
rect 5398 114438 5400 114490
rect 5344 114436 5400 114438
rect 4476 113706 4532 113708
rect 4476 113654 4478 113706
rect 4478 113654 4530 113706
rect 4530 113654 4532 113706
rect 4476 113652 4532 113654
rect 4580 113706 4636 113708
rect 4580 113654 4582 113706
rect 4582 113654 4634 113706
rect 4634 113654 4636 113706
rect 4580 113652 4636 113654
rect 4684 113706 4740 113708
rect 4684 113654 4686 113706
rect 4686 113654 4738 113706
rect 4738 113654 4740 113706
rect 4684 113652 4740 113654
rect 5136 112922 5192 112924
rect 5136 112870 5138 112922
rect 5138 112870 5190 112922
rect 5190 112870 5192 112922
rect 5136 112868 5192 112870
rect 5240 112922 5296 112924
rect 5240 112870 5242 112922
rect 5242 112870 5294 112922
rect 5294 112870 5296 112922
rect 5240 112868 5296 112870
rect 5344 112922 5400 112924
rect 5344 112870 5346 112922
rect 5346 112870 5398 112922
rect 5398 112870 5400 112922
rect 5344 112868 5400 112870
rect 2828 112418 2884 112420
rect 2828 112366 2830 112418
rect 2830 112366 2882 112418
rect 2882 112366 2884 112418
rect 2828 112364 2884 112366
rect 9212 112364 9268 112420
rect 4476 112138 4532 112140
rect 4476 112086 4478 112138
rect 4478 112086 4530 112138
rect 4530 112086 4532 112138
rect 4476 112084 4532 112086
rect 4580 112138 4636 112140
rect 4580 112086 4582 112138
rect 4582 112086 4634 112138
rect 4634 112086 4636 112138
rect 4580 112084 4636 112086
rect 4684 112138 4740 112140
rect 4684 112086 4686 112138
rect 4686 112086 4738 112138
rect 4738 112086 4740 112138
rect 4684 112084 4740 112086
rect 5136 111354 5192 111356
rect 5136 111302 5138 111354
rect 5138 111302 5190 111354
rect 5190 111302 5192 111354
rect 5136 111300 5192 111302
rect 5240 111354 5296 111356
rect 5240 111302 5242 111354
rect 5242 111302 5294 111354
rect 5294 111302 5296 111354
rect 5240 111300 5296 111302
rect 5344 111354 5400 111356
rect 5344 111302 5346 111354
rect 5346 111302 5398 111354
rect 5398 111302 5400 111354
rect 5344 111300 5400 111302
rect 4476 110570 4532 110572
rect 4476 110518 4478 110570
rect 4478 110518 4530 110570
rect 4530 110518 4532 110570
rect 4476 110516 4532 110518
rect 4580 110570 4636 110572
rect 4580 110518 4582 110570
rect 4582 110518 4634 110570
rect 4634 110518 4636 110570
rect 4580 110516 4636 110518
rect 4684 110570 4740 110572
rect 4684 110518 4686 110570
rect 4686 110518 4738 110570
rect 4738 110518 4740 110570
rect 4684 110516 4740 110518
rect 5136 109786 5192 109788
rect 5136 109734 5138 109786
rect 5138 109734 5190 109786
rect 5190 109734 5192 109786
rect 5136 109732 5192 109734
rect 5240 109786 5296 109788
rect 5240 109734 5242 109786
rect 5242 109734 5294 109786
rect 5294 109734 5296 109786
rect 5240 109732 5296 109734
rect 5344 109786 5400 109788
rect 5344 109734 5346 109786
rect 5346 109734 5398 109786
rect 5398 109734 5400 109786
rect 5344 109732 5400 109734
rect 4476 109002 4532 109004
rect 4476 108950 4478 109002
rect 4478 108950 4530 109002
rect 4530 108950 4532 109002
rect 4476 108948 4532 108950
rect 4580 109002 4636 109004
rect 4580 108950 4582 109002
rect 4582 108950 4634 109002
rect 4634 108950 4636 109002
rect 4580 108948 4636 108950
rect 4684 109002 4740 109004
rect 4684 108950 4686 109002
rect 4686 108950 4738 109002
rect 4738 108950 4740 109002
rect 4684 108948 4740 108950
rect 5136 108218 5192 108220
rect 5136 108166 5138 108218
rect 5138 108166 5190 108218
rect 5190 108166 5192 108218
rect 5136 108164 5192 108166
rect 5240 108218 5296 108220
rect 5240 108166 5242 108218
rect 5242 108166 5294 108218
rect 5294 108166 5296 108218
rect 5240 108164 5296 108166
rect 5344 108218 5400 108220
rect 5344 108166 5346 108218
rect 5346 108166 5398 108218
rect 5398 108166 5400 108218
rect 5344 108164 5400 108166
rect 4476 107434 4532 107436
rect 4476 107382 4478 107434
rect 4478 107382 4530 107434
rect 4530 107382 4532 107434
rect 4476 107380 4532 107382
rect 4580 107434 4636 107436
rect 4580 107382 4582 107434
rect 4582 107382 4634 107434
rect 4634 107382 4636 107434
rect 4580 107380 4636 107382
rect 4684 107434 4740 107436
rect 4684 107382 4686 107434
rect 4686 107382 4738 107434
rect 4738 107382 4740 107434
rect 4684 107380 4740 107382
rect 5136 106650 5192 106652
rect 5136 106598 5138 106650
rect 5138 106598 5190 106650
rect 5190 106598 5192 106650
rect 5136 106596 5192 106598
rect 5240 106650 5296 106652
rect 5240 106598 5242 106650
rect 5242 106598 5294 106650
rect 5294 106598 5296 106650
rect 5240 106596 5296 106598
rect 5344 106650 5400 106652
rect 5344 106598 5346 106650
rect 5346 106598 5398 106650
rect 5398 106598 5400 106650
rect 5344 106596 5400 106598
rect 4476 105866 4532 105868
rect 4476 105814 4478 105866
rect 4478 105814 4530 105866
rect 4530 105814 4532 105866
rect 4476 105812 4532 105814
rect 4580 105866 4636 105868
rect 4580 105814 4582 105866
rect 4582 105814 4634 105866
rect 4634 105814 4636 105866
rect 4580 105812 4636 105814
rect 4684 105866 4740 105868
rect 4684 105814 4686 105866
rect 4686 105814 4738 105866
rect 4738 105814 4740 105866
rect 4684 105812 4740 105814
rect 5136 105082 5192 105084
rect 5136 105030 5138 105082
rect 5138 105030 5190 105082
rect 5190 105030 5192 105082
rect 5136 105028 5192 105030
rect 5240 105082 5296 105084
rect 5240 105030 5242 105082
rect 5242 105030 5294 105082
rect 5294 105030 5296 105082
rect 5240 105028 5296 105030
rect 5344 105082 5400 105084
rect 5344 105030 5346 105082
rect 5346 105030 5398 105082
rect 5398 105030 5400 105082
rect 5344 105028 5400 105030
rect 4476 104298 4532 104300
rect 4476 104246 4478 104298
rect 4478 104246 4530 104298
rect 4530 104246 4532 104298
rect 4476 104244 4532 104246
rect 4580 104298 4636 104300
rect 4580 104246 4582 104298
rect 4582 104246 4634 104298
rect 4634 104246 4636 104298
rect 4580 104244 4636 104246
rect 4684 104298 4740 104300
rect 4684 104246 4686 104298
rect 4686 104246 4738 104298
rect 4738 104246 4740 104298
rect 4684 104244 4740 104246
rect 5136 103514 5192 103516
rect 5136 103462 5138 103514
rect 5138 103462 5190 103514
rect 5190 103462 5192 103514
rect 5136 103460 5192 103462
rect 5240 103514 5296 103516
rect 5240 103462 5242 103514
rect 5242 103462 5294 103514
rect 5294 103462 5296 103514
rect 5240 103460 5296 103462
rect 5344 103514 5400 103516
rect 5344 103462 5346 103514
rect 5346 103462 5398 103514
rect 5398 103462 5400 103514
rect 5344 103460 5400 103462
rect 4476 102730 4532 102732
rect 4476 102678 4478 102730
rect 4478 102678 4530 102730
rect 4530 102678 4532 102730
rect 4476 102676 4532 102678
rect 4580 102730 4636 102732
rect 4580 102678 4582 102730
rect 4582 102678 4634 102730
rect 4634 102678 4636 102730
rect 4580 102676 4636 102678
rect 4684 102730 4740 102732
rect 4684 102678 4686 102730
rect 4686 102678 4738 102730
rect 4738 102678 4740 102730
rect 4684 102676 4740 102678
rect 5136 101946 5192 101948
rect 5136 101894 5138 101946
rect 5138 101894 5190 101946
rect 5190 101894 5192 101946
rect 5136 101892 5192 101894
rect 5240 101946 5296 101948
rect 5240 101894 5242 101946
rect 5242 101894 5294 101946
rect 5294 101894 5296 101946
rect 5240 101892 5296 101894
rect 5344 101946 5400 101948
rect 5344 101894 5346 101946
rect 5346 101894 5398 101946
rect 5398 101894 5400 101946
rect 5344 101892 5400 101894
rect 7532 101612 7588 101668
rect 2492 101442 2548 101444
rect 2492 101390 2494 101442
rect 2494 101390 2546 101442
rect 2546 101390 2548 101442
rect 2492 101388 2548 101390
rect 4476 101162 4532 101164
rect 4476 101110 4478 101162
rect 4478 101110 4530 101162
rect 4530 101110 4532 101162
rect 4476 101108 4532 101110
rect 4580 101162 4636 101164
rect 4580 101110 4582 101162
rect 4582 101110 4634 101162
rect 4634 101110 4636 101162
rect 4580 101108 4636 101110
rect 4684 101162 4740 101164
rect 4684 101110 4686 101162
rect 4686 101110 4738 101162
rect 4738 101110 4740 101162
rect 4684 101108 4740 101110
rect 5136 100378 5192 100380
rect 5136 100326 5138 100378
rect 5138 100326 5190 100378
rect 5190 100326 5192 100378
rect 5136 100324 5192 100326
rect 5240 100378 5296 100380
rect 5240 100326 5242 100378
rect 5242 100326 5294 100378
rect 5294 100326 5296 100378
rect 5240 100324 5296 100326
rect 5344 100378 5400 100380
rect 5344 100326 5346 100378
rect 5346 100326 5398 100378
rect 5398 100326 5400 100378
rect 5344 100324 5400 100326
rect 4476 99594 4532 99596
rect 4476 99542 4478 99594
rect 4478 99542 4530 99594
rect 4530 99542 4532 99594
rect 4476 99540 4532 99542
rect 4580 99594 4636 99596
rect 4580 99542 4582 99594
rect 4582 99542 4634 99594
rect 4634 99542 4636 99594
rect 4580 99540 4636 99542
rect 4684 99594 4740 99596
rect 4684 99542 4686 99594
rect 4686 99542 4738 99594
rect 4738 99542 4740 99594
rect 4684 99540 4740 99542
rect 5136 98810 5192 98812
rect 5136 98758 5138 98810
rect 5138 98758 5190 98810
rect 5190 98758 5192 98810
rect 5136 98756 5192 98758
rect 5240 98810 5296 98812
rect 5240 98758 5242 98810
rect 5242 98758 5294 98810
rect 5294 98758 5296 98810
rect 5240 98756 5296 98758
rect 5344 98810 5400 98812
rect 5344 98758 5346 98810
rect 5346 98758 5398 98810
rect 5398 98758 5400 98810
rect 5344 98756 5400 98758
rect 4476 98026 4532 98028
rect 4476 97974 4478 98026
rect 4478 97974 4530 98026
rect 4530 97974 4532 98026
rect 4476 97972 4532 97974
rect 4580 98026 4636 98028
rect 4580 97974 4582 98026
rect 4582 97974 4634 98026
rect 4634 97974 4636 98026
rect 4580 97972 4636 97974
rect 4684 98026 4740 98028
rect 4684 97974 4686 98026
rect 4686 97974 4738 98026
rect 4738 97974 4740 98026
rect 4684 97972 4740 97974
rect 5136 97242 5192 97244
rect 5136 97190 5138 97242
rect 5138 97190 5190 97242
rect 5190 97190 5192 97242
rect 5136 97188 5192 97190
rect 5240 97242 5296 97244
rect 5240 97190 5242 97242
rect 5242 97190 5294 97242
rect 5294 97190 5296 97242
rect 5240 97188 5296 97190
rect 5344 97242 5400 97244
rect 5344 97190 5346 97242
rect 5346 97190 5398 97242
rect 5398 97190 5400 97242
rect 5344 97188 5400 97190
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 5136 95674 5192 95676
rect 5136 95622 5138 95674
rect 5138 95622 5190 95674
rect 5190 95622 5192 95674
rect 5136 95620 5192 95622
rect 5240 95674 5296 95676
rect 5240 95622 5242 95674
rect 5242 95622 5294 95674
rect 5294 95622 5296 95674
rect 5240 95620 5296 95622
rect 5344 95674 5400 95676
rect 5344 95622 5346 95674
rect 5346 95622 5398 95674
rect 5398 95622 5400 95674
rect 5344 95620 5400 95622
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 5136 94106 5192 94108
rect 5136 94054 5138 94106
rect 5138 94054 5190 94106
rect 5190 94054 5192 94106
rect 5136 94052 5192 94054
rect 5240 94106 5296 94108
rect 5240 94054 5242 94106
rect 5242 94054 5294 94106
rect 5294 94054 5296 94106
rect 5240 94052 5296 94054
rect 5344 94106 5400 94108
rect 5344 94054 5346 94106
rect 5346 94054 5398 94106
rect 5398 94054 5400 94106
rect 5344 94052 5400 94054
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 5136 92538 5192 92540
rect 5136 92486 5138 92538
rect 5138 92486 5190 92538
rect 5190 92486 5192 92538
rect 5136 92484 5192 92486
rect 5240 92538 5296 92540
rect 5240 92486 5242 92538
rect 5242 92486 5294 92538
rect 5294 92486 5296 92538
rect 5240 92484 5296 92486
rect 5344 92538 5400 92540
rect 5344 92486 5346 92538
rect 5346 92486 5398 92538
rect 5398 92486 5400 92538
rect 5344 92484 5400 92486
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 5136 90970 5192 90972
rect 5136 90918 5138 90970
rect 5138 90918 5190 90970
rect 5190 90918 5192 90970
rect 5136 90916 5192 90918
rect 5240 90970 5296 90972
rect 5240 90918 5242 90970
rect 5242 90918 5294 90970
rect 5294 90918 5296 90970
rect 5240 90916 5296 90918
rect 5344 90970 5400 90972
rect 5344 90918 5346 90970
rect 5346 90918 5398 90970
rect 5398 90918 5400 90970
rect 5344 90916 5400 90918
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 2492 89404 2548 89460
rect 5136 89402 5192 89404
rect 5136 89350 5138 89402
rect 5138 89350 5190 89402
rect 5190 89350 5192 89402
rect 5136 89348 5192 89350
rect 5240 89402 5296 89404
rect 5240 89350 5242 89402
rect 5242 89350 5294 89402
rect 5294 89350 5296 89402
rect 5240 89348 5296 89350
rect 5344 89402 5400 89404
rect 5344 89350 5346 89402
rect 5346 89350 5398 89402
rect 5398 89350 5400 89402
rect 5344 89348 5400 89350
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 5136 87834 5192 87836
rect 5136 87782 5138 87834
rect 5138 87782 5190 87834
rect 5190 87782 5192 87834
rect 5136 87780 5192 87782
rect 5240 87834 5296 87836
rect 5240 87782 5242 87834
rect 5242 87782 5294 87834
rect 5294 87782 5296 87834
rect 5240 87780 5296 87782
rect 5344 87834 5400 87836
rect 5344 87782 5346 87834
rect 5346 87782 5398 87834
rect 5398 87782 5400 87834
rect 5344 87780 5400 87782
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 5136 86266 5192 86268
rect 5136 86214 5138 86266
rect 5138 86214 5190 86266
rect 5190 86214 5192 86266
rect 5136 86212 5192 86214
rect 5240 86266 5296 86268
rect 5240 86214 5242 86266
rect 5242 86214 5294 86266
rect 5294 86214 5296 86266
rect 5240 86212 5296 86214
rect 5344 86266 5400 86268
rect 5344 86214 5346 86266
rect 5346 86214 5398 86266
rect 5398 86214 5400 86266
rect 5344 86212 5400 86214
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 5136 84698 5192 84700
rect 5136 84646 5138 84698
rect 5138 84646 5190 84698
rect 5190 84646 5192 84698
rect 5136 84644 5192 84646
rect 5240 84698 5296 84700
rect 5240 84646 5242 84698
rect 5242 84646 5294 84698
rect 5294 84646 5296 84698
rect 5240 84644 5296 84646
rect 5344 84698 5400 84700
rect 5344 84646 5346 84698
rect 5346 84646 5398 84698
rect 5398 84646 5400 84698
rect 5344 84644 5400 84646
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 5136 83130 5192 83132
rect 5136 83078 5138 83130
rect 5138 83078 5190 83130
rect 5190 83078 5192 83130
rect 5136 83076 5192 83078
rect 5240 83130 5296 83132
rect 5240 83078 5242 83130
rect 5242 83078 5294 83130
rect 5294 83078 5296 83130
rect 5240 83076 5296 83078
rect 5344 83130 5400 83132
rect 5344 83078 5346 83130
rect 5346 83078 5398 83130
rect 5398 83078 5400 83130
rect 5344 83076 5400 83078
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 5136 81562 5192 81564
rect 5136 81510 5138 81562
rect 5138 81510 5190 81562
rect 5190 81510 5192 81562
rect 5136 81508 5192 81510
rect 5240 81562 5296 81564
rect 5240 81510 5242 81562
rect 5242 81510 5294 81562
rect 5294 81510 5296 81562
rect 5240 81508 5296 81510
rect 5344 81562 5400 81564
rect 5344 81510 5346 81562
rect 5346 81510 5398 81562
rect 5398 81510 5400 81562
rect 5344 81508 5400 81510
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 5136 79994 5192 79996
rect 5136 79942 5138 79994
rect 5138 79942 5190 79994
rect 5190 79942 5192 79994
rect 5136 79940 5192 79942
rect 5240 79994 5296 79996
rect 5240 79942 5242 79994
rect 5242 79942 5294 79994
rect 5294 79942 5296 79994
rect 5240 79940 5296 79942
rect 5344 79994 5400 79996
rect 5344 79942 5346 79994
rect 5346 79942 5398 79994
rect 5398 79942 5400 79994
rect 5344 79940 5400 79942
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 2492 78594 2548 78596
rect 2492 78542 2494 78594
rect 2494 78542 2546 78594
rect 2546 78542 2548 78594
rect 2492 78540 2548 78542
rect 5136 78426 5192 78428
rect 5136 78374 5138 78426
rect 5138 78374 5190 78426
rect 5190 78374 5192 78426
rect 5136 78372 5192 78374
rect 5240 78426 5296 78428
rect 5240 78374 5242 78426
rect 5242 78374 5294 78426
rect 5294 78374 5296 78426
rect 5240 78372 5296 78374
rect 5344 78426 5400 78428
rect 5344 78374 5346 78426
rect 5346 78374 5398 78426
rect 5398 78374 5400 78426
rect 5344 78372 5400 78374
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 5136 76858 5192 76860
rect 5136 76806 5138 76858
rect 5138 76806 5190 76858
rect 5190 76806 5192 76858
rect 5136 76804 5192 76806
rect 5240 76858 5296 76860
rect 5240 76806 5242 76858
rect 5242 76806 5294 76858
rect 5294 76806 5296 76858
rect 5240 76804 5296 76806
rect 5344 76858 5400 76860
rect 5344 76806 5346 76858
rect 5346 76806 5398 76858
rect 5398 76806 5400 76858
rect 5344 76804 5400 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 5136 75290 5192 75292
rect 5136 75238 5138 75290
rect 5138 75238 5190 75290
rect 5190 75238 5192 75290
rect 5136 75236 5192 75238
rect 5240 75290 5296 75292
rect 5240 75238 5242 75290
rect 5242 75238 5294 75290
rect 5294 75238 5296 75290
rect 5240 75236 5296 75238
rect 5344 75290 5400 75292
rect 5344 75238 5346 75290
rect 5346 75238 5398 75290
rect 5398 75238 5400 75290
rect 5344 75236 5400 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 5136 73722 5192 73724
rect 5136 73670 5138 73722
rect 5138 73670 5190 73722
rect 5190 73670 5192 73722
rect 5136 73668 5192 73670
rect 5240 73722 5296 73724
rect 5240 73670 5242 73722
rect 5242 73670 5294 73722
rect 5294 73670 5296 73722
rect 5240 73668 5296 73670
rect 5344 73722 5400 73724
rect 5344 73670 5346 73722
rect 5346 73670 5398 73722
rect 5398 73670 5400 73722
rect 5344 73668 5400 73670
rect 7532 73164 7588 73220
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 5136 72154 5192 72156
rect 5136 72102 5138 72154
rect 5138 72102 5190 72154
rect 5190 72102 5192 72154
rect 5136 72100 5192 72102
rect 5240 72154 5296 72156
rect 5240 72102 5242 72154
rect 5242 72102 5294 72154
rect 5294 72102 5296 72154
rect 5240 72100 5296 72102
rect 5344 72154 5400 72156
rect 5344 72102 5346 72154
rect 5346 72102 5398 72154
rect 5398 72102 5400 72154
rect 5344 72100 5400 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 5136 70586 5192 70588
rect 5136 70534 5138 70586
rect 5138 70534 5190 70586
rect 5190 70534 5192 70586
rect 5136 70532 5192 70534
rect 5240 70586 5296 70588
rect 5240 70534 5242 70586
rect 5242 70534 5294 70586
rect 5294 70534 5296 70586
rect 5240 70532 5296 70534
rect 5344 70586 5400 70588
rect 5344 70534 5346 70586
rect 5346 70534 5398 70586
rect 5398 70534 5400 70586
rect 5344 70532 5400 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 5136 69018 5192 69020
rect 5136 68966 5138 69018
rect 5138 68966 5190 69018
rect 5190 68966 5192 69018
rect 5136 68964 5192 68966
rect 5240 69018 5296 69020
rect 5240 68966 5242 69018
rect 5242 68966 5294 69018
rect 5294 68966 5296 69018
rect 5240 68964 5296 68966
rect 5344 69018 5400 69020
rect 5344 68966 5346 69018
rect 5346 68966 5398 69018
rect 5398 68966 5400 69018
rect 5344 68964 5400 68966
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 5136 67450 5192 67452
rect 5136 67398 5138 67450
rect 5138 67398 5190 67450
rect 5190 67398 5192 67450
rect 5136 67396 5192 67398
rect 5240 67450 5296 67452
rect 5240 67398 5242 67450
rect 5242 67398 5294 67450
rect 5294 67398 5296 67450
rect 5240 67396 5296 67398
rect 5344 67450 5400 67452
rect 5344 67398 5346 67450
rect 5346 67398 5398 67450
rect 5398 67398 5400 67450
rect 5344 67396 5400 67398
rect 2492 66556 2548 66612
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 5136 65882 5192 65884
rect 5136 65830 5138 65882
rect 5138 65830 5190 65882
rect 5190 65830 5192 65882
rect 5136 65828 5192 65830
rect 5240 65882 5296 65884
rect 5240 65830 5242 65882
rect 5242 65830 5294 65882
rect 5294 65830 5296 65882
rect 5240 65828 5296 65830
rect 5344 65882 5400 65884
rect 5344 65830 5346 65882
rect 5346 65830 5398 65882
rect 5398 65830 5400 65882
rect 5344 65828 5400 65830
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 5136 64314 5192 64316
rect 5136 64262 5138 64314
rect 5138 64262 5190 64314
rect 5190 64262 5192 64314
rect 5136 64260 5192 64262
rect 5240 64314 5296 64316
rect 5240 64262 5242 64314
rect 5242 64262 5294 64314
rect 5294 64262 5296 64314
rect 5240 64260 5296 64262
rect 5344 64314 5400 64316
rect 5344 64262 5346 64314
rect 5346 64262 5398 64314
rect 5398 64262 5400 64314
rect 5344 64260 5400 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 5136 62746 5192 62748
rect 5136 62694 5138 62746
rect 5138 62694 5190 62746
rect 5190 62694 5192 62746
rect 5136 62692 5192 62694
rect 5240 62746 5296 62748
rect 5240 62694 5242 62746
rect 5242 62694 5294 62746
rect 5294 62694 5296 62746
rect 5240 62692 5296 62694
rect 5344 62746 5400 62748
rect 5344 62694 5346 62746
rect 5346 62694 5398 62746
rect 5398 62694 5400 62746
rect 5344 62692 5400 62694
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 5136 61178 5192 61180
rect 5136 61126 5138 61178
rect 5138 61126 5190 61178
rect 5190 61126 5192 61178
rect 5136 61124 5192 61126
rect 5240 61178 5296 61180
rect 5240 61126 5242 61178
rect 5242 61126 5294 61178
rect 5294 61126 5296 61178
rect 5240 61124 5296 61126
rect 5344 61178 5400 61180
rect 5344 61126 5346 61178
rect 5346 61126 5398 61178
rect 5398 61126 5400 61178
rect 5344 61124 5400 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 5136 59610 5192 59612
rect 5136 59558 5138 59610
rect 5138 59558 5190 59610
rect 5190 59558 5192 59610
rect 5136 59556 5192 59558
rect 5240 59610 5296 59612
rect 5240 59558 5242 59610
rect 5242 59558 5294 59610
rect 5294 59558 5296 59610
rect 5240 59556 5296 59558
rect 5344 59610 5400 59612
rect 5344 59558 5346 59610
rect 5346 59558 5398 59610
rect 5398 59558 5400 59610
rect 5344 59556 5400 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 5136 58042 5192 58044
rect 5136 57990 5138 58042
rect 5138 57990 5190 58042
rect 5190 57990 5192 58042
rect 5136 57988 5192 57990
rect 5240 58042 5296 58044
rect 5240 57990 5242 58042
rect 5242 57990 5294 58042
rect 5294 57990 5296 58042
rect 5240 57988 5296 57990
rect 5344 58042 5400 58044
rect 5344 57990 5346 58042
rect 5346 57990 5398 58042
rect 5398 57990 5400 58042
rect 5344 57988 5400 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 5136 56474 5192 56476
rect 5136 56422 5138 56474
rect 5138 56422 5190 56474
rect 5190 56422 5192 56474
rect 5136 56420 5192 56422
rect 5240 56474 5296 56476
rect 5240 56422 5242 56474
rect 5242 56422 5294 56474
rect 5294 56422 5296 56474
rect 5240 56420 5296 56422
rect 5344 56474 5400 56476
rect 5344 56422 5346 56474
rect 5346 56422 5398 56474
rect 5398 56422 5400 56474
rect 5344 56420 5400 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 5136 54906 5192 54908
rect 5136 54854 5138 54906
rect 5138 54854 5190 54906
rect 5190 54854 5192 54906
rect 5136 54852 5192 54854
rect 5240 54906 5296 54908
rect 5240 54854 5242 54906
rect 5242 54854 5294 54906
rect 5294 54854 5296 54906
rect 5240 54852 5296 54854
rect 5344 54906 5400 54908
rect 5344 54854 5346 54906
rect 5346 54854 5398 54906
rect 5398 54854 5400 54906
rect 5344 54852 5400 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 5136 53338 5192 53340
rect 5136 53286 5138 53338
rect 5138 53286 5190 53338
rect 5190 53286 5192 53338
rect 5136 53284 5192 53286
rect 5240 53338 5296 53340
rect 5240 53286 5242 53338
rect 5242 53286 5294 53338
rect 5294 53286 5296 53338
rect 5240 53284 5296 53286
rect 5344 53338 5400 53340
rect 5344 53286 5346 53338
rect 5346 53286 5398 53338
rect 5398 53286 5400 53338
rect 5344 53284 5400 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 5136 51770 5192 51772
rect 5136 51718 5138 51770
rect 5138 51718 5190 51770
rect 5190 51718 5192 51770
rect 5136 51716 5192 51718
rect 5240 51770 5296 51772
rect 5240 51718 5242 51770
rect 5242 51718 5294 51770
rect 5294 51718 5296 51770
rect 5240 51716 5296 51718
rect 5344 51770 5400 51772
rect 5344 51718 5346 51770
rect 5346 51718 5398 51770
rect 5398 51718 5400 51770
rect 5344 51716 5400 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 5136 50202 5192 50204
rect 5136 50150 5138 50202
rect 5138 50150 5190 50202
rect 5190 50150 5192 50202
rect 5136 50148 5192 50150
rect 5240 50202 5296 50204
rect 5240 50150 5242 50202
rect 5242 50150 5294 50202
rect 5294 50150 5296 50202
rect 5240 50148 5296 50150
rect 5344 50202 5400 50204
rect 5344 50150 5346 50202
rect 5346 50150 5398 50202
rect 5398 50150 5400 50202
rect 5344 50148 5400 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 5136 48634 5192 48636
rect 5136 48582 5138 48634
rect 5138 48582 5190 48634
rect 5190 48582 5192 48634
rect 5136 48580 5192 48582
rect 5240 48634 5296 48636
rect 5240 48582 5242 48634
rect 5242 48582 5294 48634
rect 5294 48582 5296 48634
rect 5240 48580 5296 48582
rect 5344 48634 5400 48636
rect 5344 48582 5346 48634
rect 5346 48582 5398 48634
rect 5398 48582 5400 48634
rect 5344 48580 5400 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 5136 47066 5192 47068
rect 5136 47014 5138 47066
rect 5138 47014 5190 47066
rect 5190 47014 5192 47066
rect 5136 47012 5192 47014
rect 5240 47066 5296 47068
rect 5240 47014 5242 47066
rect 5242 47014 5294 47066
rect 5294 47014 5296 47066
rect 5240 47012 5296 47014
rect 5344 47066 5400 47068
rect 5344 47014 5346 47066
rect 5346 47014 5398 47066
rect 5398 47014 5400 47066
rect 5344 47012 5400 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 5136 45498 5192 45500
rect 5136 45446 5138 45498
rect 5138 45446 5190 45498
rect 5190 45446 5192 45498
rect 5136 45444 5192 45446
rect 5240 45498 5296 45500
rect 5240 45446 5242 45498
rect 5242 45446 5294 45498
rect 5294 45446 5296 45498
rect 5240 45444 5296 45446
rect 5344 45498 5400 45500
rect 5344 45446 5346 45498
rect 5346 45446 5398 45498
rect 5398 45446 5400 45498
rect 5344 45444 5400 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 5136 43930 5192 43932
rect 5136 43878 5138 43930
rect 5138 43878 5190 43930
rect 5190 43878 5192 43930
rect 5136 43876 5192 43878
rect 5240 43930 5296 43932
rect 5240 43878 5242 43930
rect 5242 43878 5294 43930
rect 5294 43878 5296 43930
rect 5240 43876 5296 43878
rect 5344 43930 5400 43932
rect 5344 43878 5346 43930
rect 5346 43878 5398 43930
rect 5398 43878 5400 43930
rect 5344 43876 5400 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5136 42362 5192 42364
rect 5136 42310 5138 42362
rect 5138 42310 5190 42362
rect 5190 42310 5192 42362
rect 5136 42308 5192 42310
rect 5240 42362 5296 42364
rect 5240 42310 5242 42362
rect 5242 42310 5294 42362
rect 5294 42310 5296 42362
rect 5240 42308 5296 42310
rect 5344 42362 5400 42364
rect 5344 42310 5346 42362
rect 5346 42310 5398 42362
rect 5398 42310 5400 42362
rect 5344 42308 5400 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5136 40794 5192 40796
rect 5136 40742 5138 40794
rect 5138 40742 5190 40794
rect 5190 40742 5192 40794
rect 5136 40740 5192 40742
rect 5240 40794 5296 40796
rect 5240 40742 5242 40794
rect 5242 40742 5294 40794
rect 5294 40742 5296 40794
rect 5240 40740 5296 40742
rect 5344 40794 5400 40796
rect 5344 40742 5346 40794
rect 5346 40742 5398 40794
rect 5398 40742 5400 40794
rect 5344 40740 5400 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5136 39226 5192 39228
rect 5136 39174 5138 39226
rect 5138 39174 5190 39226
rect 5190 39174 5192 39226
rect 5136 39172 5192 39174
rect 5240 39226 5296 39228
rect 5240 39174 5242 39226
rect 5242 39174 5294 39226
rect 5294 39174 5296 39226
rect 5240 39172 5296 39174
rect 5344 39226 5400 39228
rect 5344 39174 5346 39226
rect 5346 39174 5398 39226
rect 5398 39174 5400 39226
rect 5344 39172 5400 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5136 37658 5192 37660
rect 5136 37606 5138 37658
rect 5138 37606 5190 37658
rect 5190 37606 5192 37658
rect 5136 37604 5192 37606
rect 5240 37658 5296 37660
rect 5240 37606 5242 37658
rect 5242 37606 5294 37658
rect 5294 37606 5296 37658
rect 5240 37604 5296 37606
rect 5344 37658 5400 37660
rect 5344 37606 5346 37658
rect 5346 37606 5398 37658
rect 5398 37606 5400 37658
rect 5344 37604 5400 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5136 36090 5192 36092
rect 5136 36038 5138 36090
rect 5138 36038 5190 36090
rect 5190 36038 5192 36090
rect 5136 36036 5192 36038
rect 5240 36090 5296 36092
rect 5240 36038 5242 36090
rect 5242 36038 5294 36090
rect 5294 36038 5296 36090
rect 5240 36036 5296 36038
rect 5344 36090 5400 36092
rect 5344 36038 5346 36090
rect 5346 36038 5398 36090
rect 5398 36038 5400 36090
rect 5344 36036 5400 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5136 34522 5192 34524
rect 5136 34470 5138 34522
rect 5138 34470 5190 34522
rect 5190 34470 5192 34522
rect 5136 34468 5192 34470
rect 5240 34522 5296 34524
rect 5240 34470 5242 34522
rect 5242 34470 5294 34522
rect 5294 34470 5296 34522
rect 5240 34468 5296 34470
rect 5344 34522 5400 34524
rect 5344 34470 5346 34522
rect 5346 34470 5398 34522
rect 5398 34470 5400 34522
rect 5344 34468 5400 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5136 32954 5192 32956
rect 5136 32902 5138 32954
rect 5138 32902 5190 32954
rect 5190 32902 5192 32954
rect 5136 32900 5192 32902
rect 5240 32954 5296 32956
rect 5240 32902 5242 32954
rect 5242 32902 5294 32954
rect 5294 32902 5296 32954
rect 5240 32900 5296 32902
rect 5344 32954 5400 32956
rect 5344 32902 5346 32954
rect 5346 32902 5398 32954
rect 5398 32902 5400 32954
rect 5344 32900 5400 32902
rect 2492 32284 2548 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5136 31386 5192 31388
rect 5136 31334 5138 31386
rect 5138 31334 5190 31386
rect 5190 31334 5192 31386
rect 5136 31332 5192 31334
rect 5240 31386 5296 31388
rect 5240 31334 5242 31386
rect 5242 31334 5294 31386
rect 5294 31334 5296 31386
rect 5240 31332 5296 31334
rect 5344 31386 5400 31388
rect 5344 31334 5346 31386
rect 5346 31334 5398 31386
rect 5398 31334 5400 31386
rect 5344 31332 5400 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5136 29818 5192 29820
rect 5136 29766 5138 29818
rect 5138 29766 5190 29818
rect 5190 29766 5192 29818
rect 5136 29764 5192 29766
rect 5240 29818 5296 29820
rect 5240 29766 5242 29818
rect 5242 29766 5294 29818
rect 5294 29766 5296 29818
rect 5240 29764 5296 29766
rect 5344 29818 5400 29820
rect 5344 29766 5346 29818
rect 5346 29766 5398 29818
rect 5398 29766 5400 29818
rect 5344 29764 5400 29766
rect 2380 29372 2436 29428
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 5136 28250 5192 28252
rect 5136 28198 5138 28250
rect 5138 28198 5190 28250
rect 5190 28198 5192 28250
rect 5136 28196 5192 28198
rect 5240 28250 5296 28252
rect 5240 28198 5242 28250
rect 5242 28198 5294 28250
rect 5294 28198 5296 28250
rect 5240 28196 5296 28198
rect 5344 28250 5400 28252
rect 5344 28198 5346 28250
rect 5346 28198 5398 28250
rect 5398 28198 5400 28250
rect 5344 28196 5400 28198
rect 9212 27692 9268 27748
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5136 26682 5192 26684
rect 5136 26630 5138 26682
rect 5138 26630 5190 26682
rect 5190 26630 5192 26682
rect 5136 26628 5192 26630
rect 5240 26682 5296 26684
rect 5240 26630 5242 26682
rect 5242 26630 5294 26682
rect 5294 26630 5296 26682
rect 5240 26628 5296 26630
rect 5344 26682 5400 26684
rect 5344 26630 5346 26682
rect 5346 26630 5398 26682
rect 5398 26630 5400 26682
rect 5344 26628 5400 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5136 25114 5192 25116
rect 5136 25062 5138 25114
rect 5138 25062 5190 25114
rect 5190 25062 5192 25114
rect 5136 25060 5192 25062
rect 5240 25114 5296 25116
rect 5240 25062 5242 25114
rect 5242 25062 5294 25114
rect 5294 25062 5296 25114
rect 5240 25060 5296 25062
rect 5344 25114 5400 25116
rect 5344 25062 5346 25114
rect 5346 25062 5398 25114
rect 5398 25062 5400 25114
rect 5344 25060 5400 25062
rect 17724 135100 17780 135156
rect 14252 78540 14308 78596
rect 17612 78594 17668 78596
rect 17612 78542 17614 78594
rect 17614 78542 17666 78594
rect 17666 78542 17668 78594
rect 17612 78540 17668 78542
rect 15932 76524 15988 76580
rect 17612 76524 17668 76580
rect 17612 76354 17668 76356
rect 17612 76302 17614 76354
rect 17614 76302 17666 76354
rect 17666 76302 17668 76354
rect 17612 76300 17668 76302
rect 17500 75682 17556 75684
rect 17500 75630 17502 75682
rect 17502 75630 17554 75682
rect 17554 75630 17556 75682
rect 17500 75628 17556 75630
rect 17500 74786 17556 74788
rect 17500 74734 17502 74786
rect 17502 74734 17554 74786
rect 17554 74734 17556 74786
rect 17500 74732 17556 74734
rect 17500 73218 17556 73220
rect 17500 73166 17502 73218
rect 17502 73166 17554 73218
rect 17554 73166 17556 73218
rect 17500 73164 17556 73166
rect 15932 55244 15988 55300
rect 14252 44268 14308 44324
rect 17612 36258 17668 36260
rect 17612 36206 17614 36258
rect 17614 36206 17666 36258
rect 17666 36206 17668 36258
rect 17612 36204 17668 36206
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 12572 24332 12628 24388
rect 12684 35532 12740 35588
rect 4684 24276 4740 24278
rect 5136 23546 5192 23548
rect 5136 23494 5138 23546
rect 5138 23494 5190 23546
rect 5190 23494 5192 23546
rect 5136 23492 5192 23494
rect 5240 23546 5296 23548
rect 5240 23494 5242 23546
rect 5242 23494 5294 23546
rect 5294 23494 5296 23546
rect 5240 23492 5296 23494
rect 5344 23546 5400 23548
rect 5344 23494 5346 23546
rect 5346 23494 5398 23546
rect 5398 23494 5400 23546
rect 5344 23492 5400 23494
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5136 21978 5192 21980
rect 5136 21926 5138 21978
rect 5138 21926 5190 21978
rect 5190 21926 5192 21978
rect 5136 21924 5192 21926
rect 5240 21978 5296 21980
rect 5240 21926 5242 21978
rect 5242 21926 5294 21978
rect 5294 21926 5296 21978
rect 5240 21924 5296 21926
rect 5344 21978 5400 21980
rect 5344 21926 5346 21978
rect 5346 21926 5398 21978
rect 5398 21926 5400 21978
rect 5344 21924 5400 21926
rect 1708 21420 1764 21476
rect 2492 21474 2548 21476
rect 2492 21422 2494 21474
rect 2494 21422 2546 21474
rect 2546 21422 2548 21474
rect 2492 21420 2548 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1708 20860 1764 20916
rect 5136 20410 5192 20412
rect 5136 20358 5138 20410
rect 5138 20358 5190 20410
rect 5190 20358 5192 20410
rect 5136 20356 5192 20358
rect 5240 20410 5296 20412
rect 5240 20358 5242 20410
rect 5242 20358 5294 20410
rect 5294 20358 5296 20410
rect 5240 20356 5296 20358
rect 5344 20410 5400 20412
rect 5344 20358 5346 20410
rect 5346 20358 5398 20410
rect 5398 20358 5400 20410
rect 5344 20356 5400 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5136 18842 5192 18844
rect 5136 18790 5138 18842
rect 5138 18790 5190 18842
rect 5190 18790 5192 18842
rect 5136 18788 5192 18790
rect 5240 18842 5296 18844
rect 5240 18790 5242 18842
rect 5242 18790 5294 18842
rect 5294 18790 5296 18842
rect 5240 18788 5296 18790
rect 5344 18842 5400 18844
rect 5344 18790 5346 18842
rect 5346 18790 5398 18842
rect 5398 18790 5400 18842
rect 5344 18788 5400 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5136 17274 5192 17276
rect 5136 17222 5138 17274
rect 5138 17222 5190 17274
rect 5190 17222 5192 17274
rect 5136 17220 5192 17222
rect 5240 17274 5296 17276
rect 5240 17222 5242 17274
rect 5242 17222 5294 17274
rect 5294 17222 5296 17274
rect 5240 17220 5296 17222
rect 5344 17274 5400 17276
rect 5344 17222 5346 17274
rect 5346 17222 5398 17274
rect 5398 17222 5400 17274
rect 5344 17220 5400 17222
rect 1708 17052 1764 17108
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 5136 15706 5192 15708
rect 5136 15654 5138 15706
rect 5138 15654 5190 15706
rect 5190 15654 5192 15706
rect 5136 15652 5192 15654
rect 5240 15706 5296 15708
rect 5240 15654 5242 15706
rect 5242 15654 5294 15706
rect 5294 15654 5296 15706
rect 5240 15652 5296 15654
rect 5344 15706 5400 15708
rect 5344 15654 5346 15706
rect 5346 15654 5398 15706
rect 5398 15654 5400 15706
rect 5344 15652 5400 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5136 14138 5192 14140
rect 5136 14086 5138 14138
rect 5138 14086 5190 14138
rect 5190 14086 5192 14138
rect 5136 14084 5192 14086
rect 5240 14138 5296 14140
rect 5240 14086 5242 14138
rect 5242 14086 5294 14138
rect 5294 14086 5296 14138
rect 5240 14084 5296 14086
rect 5344 14138 5400 14140
rect 5344 14086 5346 14138
rect 5346 14086 5398 14138
rect 5398 14086 5400 14138
rect 5344 14084 5400 14086
rect 1708 13244 1764 13300
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5136 12570 5192 12572
rect 5136 12518 5138 12570
rect 5138 12518 5190 12570
rect 5190 12518 5192 12570
rect 5136 12516 5192 12518
rect 5240 12570 5296 12572
rect 5240 12518 5242 12570
rect 5242 12518 5294 12570
rect 5294 12518 5296 12570
rect 5240 12516 5296 12518
rect 5344 12570 5400 12572
rect 5344 12518 5346 12570
rect 5346 12518 5398 12570
rect 5398 12518 5400 12570
rect 5344 12516 5400 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5136 11002 5192 11004
rect 5136 10950 5138 11002
rect 5138 10950 5190 11002
rect 5190 10950 5192 11002
rect 5136 10948 5192 10950
rect 5240 11002 5296 11004
rect 5240 10950 5242 11002
rect 5242 10950 5294 11002
rect 5294 10950 5296 11002
rect 5240 10948 5296 10950
rect 5344 11002 5400 11004
rect 5344 10950 5346 11002
rect 5346 10950 5398 11002
rect 5398 10950 5400 11002
rect 5344 10948 5400 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2044 9602 2100 9604
rect 2044 9550 2046 9602
rect 2046 9550 2098 9602
rect 2098 9550 2100 9602
rect 2044 9548 2100 9550
rect 1708 9436 1764 9492
rect 17612 35586 17668 35588
rect 17612 35534 17614 35586
rect 17614 35534 17666 35586
rect 17666 35534 17668 35586
rect 17612 35532 17668 35534
rect 16940 34636 16996 34692
rect 17724 20412 17780 20468
rect 35856 156826 35912 156828
rect 35856 156774 35858 156826
rect 35858 156774 35910 156826
rect 35910 156774 35912 156826
rect 35856 156772 35912 156774
rect 35960 156826 36016 156828
rect 35960 156774 35962 156826
rect 35962 156774 36014 156826
rect 36014 156774 36016 156826
rect 35960 156772 36016 156774
rect 36064 156826 36120 156828
rect 36064 156774 36066 156826
rect 36066 156774 36118 156826
rect 36118 156774 36120 156826
rect 36064 156772 36120 156774
rect 41916 156604 41972 156660
rect 43708 156658 43764 156660
rect 43708 156606 43710 156658
rect 43710 156606 43762 156658
rect 43762 156606 43764 156658
rect 43708 156604 43764 156606
rect 42812 156322 42868 156324
rect 42812 156270 42814 156322
rect 42814 156270 42866 156322
rect 42866 156270 42868 156322
rect 42812 156268 42868 156270
rect 66576 156826 66632 156828
rect 66576 156774 66578 156826
rect 66578 156774 66630 156826
rect 66630 156774 66632 156826
rect 66576 156772 66632 156774
rect 66680 156826 66736 156828
rect 66680 156774 66682 156826
rect 66682 156774 66734 156826
rect 66734 156774 66736 156826
rect 66680 156772 66736 156774
rect 66784 156826 66840 156828
rect 66784 156774 66786 156826
rect 66786 156774 66838 156826
rect 66838 156774 66840 156826
rect 66784 156772 66840 156774
rect 64764 156604 64820 156660
rect 63756 156492 63812 156548
rect 56252 156268 56308 156324
rect 35196 156042 35252 156044
rect 35196 155990 35198 156042
rect 35198 155990 35250 156042
rect 35250 155990 35252 156042
rect 35196 155988 35252 155990
rect 35300 156042 35356 156044
rect 35300 155990 35302 156042
rect 35302 155990 35354 156042
rect 35354 155990 35356 156042
rect 35300 155988 35356 155990
rect 35404 156042 35460 156044
rect 35404 155990 35406 156042
rect 35406 155990 35458 156042
rect 35458 155990 35460 156042
rect 35404 155988 35460 155990
rect 35856 155258 35912 155260
rect 35856 155206 35858 155258
rect 35858 155206 35910 155258
rect 35910 155206 35912 155258
rect 35856 155204 35912 155206
rect 35960 155258 36016 155260
rect 35960 155206 35962 155258
rect 35962 155206 36014 155258
rect 36014 155206 36016 155258
rect 35960 155204 36016 155206
rect 36064 155258 36120 155260
rect 36064 155206 36066 155258
rect 36066 155206 36118 155258
rect 36118 155206 36120 155258
rect 36064 155204 36120 155206
rect 35196 154474 35252 154476
rect 35196 154422 35198 154474
rect 35198 154422 35250 154474
rect 35250 154422 35252 154474
rect 35196 154420 35252 154422
rect 35300 154474 35356 154476
rect 35300 154422 35302 154474
rect 35302 154422 35354 154474
rect 35354 154422 35356 154474
rect 35300 154420 35356 154422
rect 35404 154474 35460 154476
rect 35404 154422 35406 154474
rect 35406 154422 35458 154474
rect 35458 154422 35460 154474
rect 35404 154420 35460 154422
rect 35856 153690 35912 153692
rect 35856 153638 35858 153690
rect 35858 153638 35910 153690
rect 35910 153638 35912 153690
rect 35856 153636 35912 153638
rect 35960 153690 36016 153692
rect 35960 153638 35962 153690
rect 35962 153638 36014 153690
rect 36014 153638 36016 153690
rect 35960 153636 36016 153638
rect 36064 153690 36120 153692
rect 36064 153638 36066 153690
rect 36066 153638 36118 153690
rect 36118 153638 36120 153690
rect 36064 153636 36120 153638
rect 35196 152906 35252 152908
rect 35196 152854 35198 152906
rect 35198 152854 35250 152906
rect 35250 152854 35252 152906
rect 35196 152852 35252 152854
rect 35300 152906 35356 152908
rect 35300 152854 35302 152906
rect 35302 152854 35354 152906
rect 35354 152854 35356 152906
rect 35300 152852 35356 152854
rect 35404 152906 35460 152908
rect 35404 152854 35406 152906
rect 35406 152854 35458 152906
rect 35458 152854 35460 152906
rect 35404 152852 35460 152854
rect 35856 152122 35912 152124
rect 35856 152070 35858 152122
rect 35858 152070 35910 152122
rect 35910 152070 35912 152122
rect 35856 152068 35912 152070
rect 35960 152122 36016 152124
rect 35960 152070 35962 152122
rect 35962 152070 36014 152122
rect 36014 152070 36016 152122
rect 35960 152068 36016 152070
rect 36064 152122 36120 152124
rect 36064 152070 36066 152122
rect 36066 152070 36118 152122
rect 36118 152070 36120 152122
rect 36064 152068 36120 152070
rect 35196 151338 35252 151340
rect 35196 151286 35198 151338
rect 35198 151286 35250 151338
rect 35250 151286 35252 151338
rect 35196 151284 35252 151286
rect 35300 151338 35356 151340
rect 35300 151286 35302 151338
rect 35302 151286 35354 151338
rect 35354 151286 35356 151338
rect 35300 151284 35356 151286
rect 35404 151338 35460 151340
rect 35404 151286 35406 151338
rect 35406 151286 35458 151338
rect 35458 151286 35460 151338
rect 35404 151284 35460 151286
rect 35856 150554 35912 150556
rect 35856 150502 35858 150554
rect 35858 150502 35910 150554
rect 35910 150502 35912 150554
rect 35856 150500 35912 150502
rect 35960 150554 36016 150556
rect 35960 150502 35962 150554
rect 35962 150502 36014 150554
rect 36014 150502 36016 150554
rect 35960 150500 36016 150502
rect 36064 150554 36120 150556
rect 36064 150502 36066 150554
rect 36066 150502 36118 150554
rect 36118 150502 36120 150554
rect 36064 150500 36120 150502
rect 35196 149770 35252 149772
rect 35196 149718 35198 149770
rect 35198 149718 35250 149770
rect 35250 149718 35252 149770
rect 35196 149716 35252 149718
rect 35300 149770 35356 149772
rect 35300 149718 35302 149770
rect 35302 149718 35354 149770
rect 35354 149718 35356 149770
rect 35300 149716 35356 149718
rect 35404 149770 35460 149772
rect 35404 149718 35406 149770
rect 35406 149718 35458 149770
rect 35458 149718 35460 149770
rect 35404 149716 35460 149718
rect 35856 148986 35912 148988
rect 35856 148934 35858 148986
rect 35858 148934 35910 148986
rect 35910 148934 35912 148986
rect 35856 148932 35912 148934
rect 35960 148986 36016 148988
rect 35960 148934 35962 148986
rect 35962 148934 36014 148986
rect 36014 148934 36016 148986
rect 35960 148932 36016 148934
rect 36064 148986 36120 148988
rect 36064 148934 36066 148986
rect 36066 148934 36118 148986
rect 36118 148934 36120 148986
rect 36064 148932 36120 148934
rect 35196 148202 35252 148204
rect 35196 148150 35198 148202
rect 35198 148150 35250 148202
rect 35250 148150 35252 148202
rect 35196 148148 35252 148150
rect 35300 148202 35356 148204
rect 35300 148150 35302 148202
rect 35302 148150 35354 148202
rect 35354 148150 35356 148202
rect 35300 148148 35356 148150
rect 35404 148202 35460 148204
rect 35404 148150 35406 148202
rect 35406 148150 35458 148202
rect 35458 148150 35460 148202
rect 35404 148148 35460 148150
rect 35856 147418 35912 147420
rect 35856 147366 35858 147418
rect 35858 147366 35910 147418
rect 35910 147366 35912 147418
rect 35856 147364 35912 147366
rect 35960 147418 36016 147420
rect 35960 147366 35962 147418
rect 35962 147366 36014 147418
rect 36014 147366 36016 147418
rect 35960 147364 36016 147366
rect 36064 147418 36120 147420
rect 36064 147366 36066 147418
rect 36066 147366 36118 147418
rect 36118 147366 36120 147418
rect 36064 147364 36120 147366
rect 35196 146634 35252 146636
rect 35196 146582 35198 146634
rect 35198 146582 35250 146634
rect 35250 146582 35252 146634
rect 35196 146580 35252 146582
rect 35300 146634 35356 146636
rect 35300 146582 35302 146634
rect 35302 146582 35354 146634
rect 35354 146582 35356 146634
rect 35300 146580 35356 146582
rect 35404 146634 35460 146636
rect 35404 146582 35406 146634
rect 35406 146582 35458 146634
rect 35458 146582 35460 146634
rect 35404 146580 35460 146582
rect 35856 145850 35912 145852
rect 35856 145798 35858 145850
rect 35858 145798 35910 145850
rect 35910 145798 35912 145850
rect 35856 145796 35912 145798
rect 35960 145850 36016 145852
rect 35960 145798 35962 145850
rect 35962 145798 36014 145850
rect 36014 145798 36016 145850
rect 35960 145796 36016 145798
rect 36064 145850 36120 145852
rect 36064 145798 36066 145850
rect 36066 145798 36118 145850
rect 36118 145798 36120 145850
rect 36064 145796 36120 145798
rect 35196 145066 35252 145068
rect 35196 145014 35198 145066
rect 35198 145014 35250 145066
rect 35250 145014 35252 145066
rect 35196 145012 35252 145014
rect 35300 145066 35356 145068
rect 35300 145014 35302 145066
rect 35302 145014 35354 145066
rect 35354 145014 35356 145066
rect 35300 145012 35356 145014
rect 35404 145066 35460 145068
rect 35404 145014 35406 145066
rect 35406 145014 35458 145066
rect 35458 145014 35460 145066
rect 35404 145012 35460 145014
rect 26012 124124 26068 124180
rect 56252 41132 56308 41188
rect 66556 156658 66612 156660
rect 66556 156606 66558 156658
rect 66558 156606 66610 156658
rect 66610 156606 66612 156658
rect 66556 156604 66612 156606
rect 65100 156380 65156 156436
rect 64428 156268 64484 156324
rect 64428 41244 64484 41300
rect 63756 41020 63812 41076
rect 61740 38108 61796 38164
rect 26012 37996 26068 38052
rect 51436 37996 51492 38052
rect 44156 24332 44212 24388
rect 59052 37996 59108 38052
rect 53900 27692 53956 27748
rect 51436 22316 51492 22372
rect 44156 21756 44212 21812
rect 22764 18396 22820 18452
rect 44716 21196 44772 21252
rect 35856 17274 35912 17276
rect 35856 17222 35858 17274
rect 35858 17222 35910 17274
rect 35910 17222 35912 17274
rect 35856 17220 35912 17222
rect 35960 17274 36016 17276
rect 35960 17222 35962 17274
rect 35962 17222 36014 17274
rect 36014 17222 36016 17274
rect 35960 17220 36016 17222
rect 36064 17274 36120 17276
rect 36064 17222 36066 17274
rect 36066 17222 36118 17274
rect 36118 17222 36120 17274
rect 36064 17220 36120 17222
rect 48300 20412 48356 20468
rect 53900 21756 53956 21812
rect 55132 21644 55188 21700
rect 61740 22316 61796 22372
rect 65324 156322 65380 156324
rect 65324 156270 65326 156322
rect 65326 156270 65378 156322
rect 65378 156270 65380 156322
rect 65324 156268 65380 156270
rect 87612 156546 87668 156548
rect 87612 156494 87614 156546
rect 87614 156494 87666 156546
rect 87666 156494 87668 156546
rect 87612 156492 87668 156494
rect 97296 156826 97352 156828
rect 97296 156774 97298 156826
rect 97298 156774 97350 156826
rect 97350 156774 97352 156826
rect 97296 156772 97352 156774
rect 97400 156826 97456 156828
rect 97400 156774 97402 156826
rect 97402 156774 97454 156826
rect 97454 156774 97456 156826
rect 97400 156772 97456 156774
rect 97504 156826 97560 156828
rect 97504 156774 97506 156826
rect 97506 156774 97558 156826
rect 97558 156774 97560 156826
rect 97504 156772 97560 156774
rect 111132 156322 111188 156324
rect 111132 156270 111134 156322
rect 111134 156270 111186 156322
rect 111186 156270 111188 156322
rect 111132 156268 111188 156270
rect 128016 156826 128072 156828
rect 128016 156774 128018 156826
rect 128018 156774 128070 156826
rect 128070 156774 128072 156826
rect 128016 156772 128072 156774
rect 128120 156826 128176 156828
rect 128120 156774 128122 156826
rect 128122 156774 128174 156826
rect 128174 156774 128176 156826
rect 128120 156772 128176 156774
rect 128224 156826 128280 156828
rect 128224 156774 128226 156826
rect 128226 156774 128278 156826
rect 128278 156774 128280 156826
rect 128224 156772 128280 156774
rect 134204 156604 134260 156660
rect 135100 156658 135156 156660
rect 135100 156606 135102 156658
rect 135102 156606 135154 156658
rect 135154 156606 135156 156658
rect 135100 156604 135156 156606
rect 65916 156042 65972 156044
rect 65916 155990 65918 156042
rect 65918 155990 65970 156042
rect 65970 155990 65972 156042
rect 65916 155988 65972 155990
rect 66020 156042 66076 156044
rect 66020 155990 66022 156042
rect 66022 155990 66074 156042
rect 66074 155990 66076 156042
rect 66020 155988 66076 155990
rect 66124 156042 66180 156044
rect 66124 155990 66126 156042
rect 66126 155990 66178 156042
rect 66178 155990 66180 156042
rect 66124 155988 66180 155990
rect 96636 156042 96692 156044
rect 96636 155990 96638 156042
rect 96638 155990 96690 156042
rect 96690 155990 96692 156042
rect 96636 155988 96692 155990
rect 96740 156042 96796 156044
rect 96740 155990 96742 156042
rect 96742 155990 96794 156042
rect 96794 155990 96796 156042
rect 96740 155988 96796 155990
rect 96844 156042 96900 156044
rect 96844 155990 96846 156042
rect 96846 155990 96898 156042
rect 96898 155990 96900 156042
rect 96844 155988 96900 155990
rect 127356 156042 127412 156044
rect 127356 155990 127358 156042
rect 127358 155990 127410 156042
rect 127410 155990 127412 156042
rect 127356 155988 127412 155990
rect 127460 156042 127516 156044
rect 127460 155990 127462 156042
rect 127462 155990 127514 156042
rect 127514 155990 127516 156042
rect 127460 155988 127516 155990
rect 127564 156042 127620 156044
rect 127564 155990 127566 156042
rect 127566 155990 127618 156042
rect 127618 155990 127620 156042
rect 127564 155988 127620 155990
rect 66576 155258 66632 155260
rect 66576 155206 66578 155258
rect 66578 155206 66630 155258
rect 66630 155206 66632 155258
rect 66576 155204 66632 155206
rect 66680 155258 66736 155260
rect 66680 155206 66682 155258
rect 66682 155206 66734 155258
rect 66734 155206 66736 155258
rect 66680 155204 66736 155206
rect 66784 155258 66840 155260
rect 66784 155206 66786 155258
rect 66786 155206 66838 155258
rect 66838 155206 66840 155258
rect 66784 155204 66840 155206
rect 97296 155258 97352 155260
rect 97296 155206 97298 155258
rect 97298 155206 97350 155258
rect 97350 155206 97352 155258
rect 97296 155204 97352 155206
rect 97400 155258 97456 155260
rect 97400 155206 97402 155258
rect 97402 155206 97454 155258
rect 97454 155206 97456 155258
rect 97400 155204 97456 155206
rect 97504 155258 97560 155260
rect 97504 155206 97506 155258
rect 97506 155206 97558 155258
rect 97558 155206 97560 155258
rect 97504 155204 97560 155206
rect 128016 155258 128072 155260
rect 128016 155206 128018 155258
rect 128018 155206 128070 155258
rect 128070 155206 128072 155258
rect 128016 155204 128072 155206
rect 128120 155258 128176 155260
rect 128120 155206 128122 155258
rect 128122 155206 128174 155258
rect 128174 155206 128176 155258
rect 128120 155204 128176 155206
rect 128224 155258 128280 155260
rect 128224 155206 128226 155258
rect 128226 155206 128278 155258
rect 128278 155206 128280 155258
rect 128224 155204 128280 155206
rect 65916 154474 65972 154476
rect 65916 154422 65918 154474
rect 65918 154422 65970 154474
rect 65970 154422 65972 154474
rect 65916 154420 65972 154422
rect 66020 154474 66076 154476
rect 66020 154422 66022 154474
rect 66022 154422 66074 154474
rect 66074 154422 66076 154474
rect 66020 154420 66076 154422
rect 66124 154474 66180 154476
rect 66124 154422 66126 154474
rect 66126 154422 66178 154474
rect 66178 154422 66180 154474
rect 66124 154420 66180 154422
rect 96636 154474 96692 154476
rect 96636 154422 96638 154474
rect 96638 154422 96690 154474
rect 96690 154422 96692 154474
rect 96636 154420 96692 154422
rect 96740 154474 96796 154476
rect 96740 154422 96742 154474
rect 96742 154422 96794 154474
rect 96794 154422 96796 154474
rect 96740 154420 96796 154422
rect 96844 154474 96900 154476
rect 96844 154422 96846 154474
rect 96846 154422 96898 154474
rect 96898 154422 96900 154474
rect 96844 154420 96900 154422
rect 127356 154474 127412 154476
rect 127356 154422 127358 154474
rect 127358 154422 127410 154474
rect 127410 154422 127412 154474
rect 127356 154420 127412 154422
rect 127460 154474 127516 154476
rect 127460 154422 127462 154474
rect 127462 154422 127514 154474
rect 127514 154422 127516 154474
rect 127460 154420 127516 154422
rect 127564 154474 127620 154476
rect 127564 154422 127566 154474
rect 127566 154422 127618 154474
rect 127618 154422 127620 154474
rect 127564 154420 127620 154422
rect 66576 153690 66632 153692
rect 66576 153638 66578 153690
rect 66578 153638 66630 153690
rect 66630 153638 66632 153690
rect 66576 153636 66632 153638
rect 66680 153690 66736 153692
rect 66680 153638 66682 153690
rect 66682 153638 66734 153690
rect 66734 153638 66736 153690
rect 66680 153636 66736 153638
rect 66784 153690 66840 153692
rect 66784 153638 66786 153690
rect 66786 153638 66838 153690
rect 66838 153638 66840 153690
rect 66784 153636 66840 153638
rect 97296 153690 97352 153692
rect 97296 153638 97298 153690
rect 97298 153638 97350 153690
rect 97350 153638 97352 153690
rect 97296 153636 97352 153638
rect 97400 153690 97456 153692
rect 97400 153638 97402 153690
rect 97402 153638 97454 153690
rect 97454 153638 97456 153690
rect 97400 153636 97456 153638
rect 97504 153690 97560 153692
rect 97504 153638 97506 153690
rect 97506 153638 97558 153690
rect 97558 153638 97560 153690
rect 97504 153636 97560 153638
rect 128016 153690 128072 153692
rect 128016 153638 128018 153690
rect 128018 153638 128070 153690
rect 128070 153638 128072 153690
rect 128016 153636 128072 153638
rect 128120 153690 128176 153692
rect 128120 153638 128122 153690
rect 128122 153638 128174 153690
rect 128174 153638 128176 153690
rect 128120 153636 128176 153638
rect 128224 153690 128280 153692
rect 128224 153638 128226 153690
rect 128226 153638 128278 153690
rect 128278 153638 128280 153690
rect 128224 153636 128280 153638
rect 65916 152906 65972 152908
rect 65916 152854 65918 152906
rect 65918 152854 65970 152906
rect 65970 152854 65972 152906
rect 65916 152852 65972 152854
rect 66020 152906 66076 152908
rect 66020 152854 66022 152906
rect 66022 152854 66074 152906
rect 66074 152854 66076 152906
rect 66020 152852 66076 152854
rect 66124 152906 66180 152908
rect 66124 152854 66126 152906
rect 66126 152854 66178 152906
rect 66178 152854 66180 152906
rect 66124 152852 66180 152854
rect 96636 152906 96692 152908
rect 96636 152854 96638 152906
rect 96638 152854 96690 152906
rect 96690 152854 96692 152906
rect 96636 152852 96692 152854
rect 96740 152906 96796 152908
rect 96740 152854 96742 152906
rect 96742 152854 96794 152906
rect 96794 152854 96796 152906
rect 96740 152852 96796 152854
rect 96844 152906 96900 152908
rect 96844 152854 96846 152906
rect 96846 152854 96898 152906
rect 96898 152854 96900 152906
rect 96844 152852 96900 152854
rect 127356 152906 127412 152908
rect 127356 152854 127358 152906
rect 127358 152854 127410 152906
rect 127410 152854 127412 152906
rect 127356 152852 127412 152854
rect 127460 152906 127516 152908
rect 127460 152854 127462 152906
rect 127462 152854 127514 152906
rect 127514 152854 127516 152906
rect 127460 152852 127516 152854
rect 127564 152906 127620 152908
rect 127564 152854 127566 152906
rect 127566 152854 127618 152906
rect 127618 152854 127620 152906
rect 127564 152852 127620 152854
rect 66576 152122 66632 152124
rect 66576 152070 66578 152122
rect 66578 152070 66630 152122
rect 66630 152070 66632 152122
rect 66576 152068 66632 152070
rect 66680 152122 66736 152124
rect 66680 152070 66682 152122
rect 66682 152070 66734 152122
rect 66734 152070 66736 152122
rect 66680 152068 66736 152070
rect 66784 152122 66840 152124
rect 66784 152070 66786 152122
rect 66786 152070 66838 152122
rect 66838 152070 66840 152122
rect 66784 152068 66840 152070
rect 97296 152122 97352 152124
rect 97296 152070 97298 152122
rect 97298 152070 97350 152122
rect 97350 152070 97352 152122
rect 97296 152068 97352 152070
rect 97400 152122 97456 152124
rect 97400 152070 97402 152122
rect 97402 152070 97454 152122
rect 97454 152070 97456 152122
rect 97400 152068 97456 152070
rect 97504 152122 97560 152124
rect 97504 152070 97506 152122
rect 97506 152070 97558 152122
rect 97558 152070 97560 152122
rect 97504 152068 97560 152070
rect 128016 152122 128072 152124
rect 128016 152070 128018 152122
rect 128018 152070 128070 152122
rect 128070 152070 128072 152122
rect 128016 152068 128072 152070
rect 128120 152122 128176 152124
rect 128120 152070 128122 152122
rect 128122 152070 128174 152122
rect 128174 152070 128176 152122
rect 128120 152068 128176 152070
rect 128224 152122 128280 152124
rect 128224 152070 128226 152122
rect 128226 152070 128278 152122
rect 128278 152070 128280 152122
rect 128224 152068 128280 152070
rect 65916 151338 65972 151340
rect 65916 151286 65918 151338
rect 65918 151286 65970 151338
rect 65970 151286 65972 151338
rect 65916 151284 65972 151286
rect 66020 151338 66076 151340
rect 66020 151286 66022 151338
rect 66022 151286 66074 151338
rect 66074 151286 66076 151338
rect 66020 151284 66076 151286
rect 66124 151338 66180 151340
rect 66124 151286 66126 151338
rect 66126 151286 66178 151338
rect 66178 151286 66180 151338
rect 66124 151284 66180 151286
rect 96636 151338 96692 151340
rect 96636 151286 96638 151338
rect 96638 151286 96690 151338
rect 96690 151286 96692 151338
rect 96636 151284 96692 151286
rect 96740 151338 96796 151340
rect 96740 151286 96742 151338
rect 96742 151286 96794 151338
rect 96794 151286 96796 151338
rect 96740 151284 96796 151286
rect 96844 151338 96900 151340
rect 96844 151286 96846 151338
rect 96846 151286 96898 151338
rect 96898 151286 96900 151338
rect 96844 151284 96900 151286
rect 127356 151338 127412 151340
rect 127356 151286 127358 151338
rect 127358 151286 127410 151338
rect 127410 151286 127412 151338
rect 127356 151284 127412 151286
rect 127460 151338 127516 151340
rect 127460 151286 127462 151338
rect 127462 151286 127514 151338
rect 127514 151286 127516 151338
rect 127460 151284 127516 151286
rect 127564 151338 127620 151340
rect 127564 151286 127566 151338
rect 127566 151286 127618 151338
rect 127618 151286 127620 151338
rect 127564 151284 127620 151286
rect 66576 150554 66632 150556
rect 66576 150502 66578 150554
rect 66578 150502 66630 150554
rect 66630 150502 66632 150554
rect 66576 150500 66632 150502
rect 66680 150554 66736 150556
rect 66680 150502 66682 150554
rect 66682 150502 66734 150554
rect 66734 150502 66736 150554
rect 66680 150500 66736 150502
rect 66784 150554 66840 150556
rect 66784 150502 66786 150554
rect 66786 150502 66838 150554
rect 66838 150502 66840 150554
rect 66784 150500 66840 150502
rect 97296 150554 97352 150556
rect 97296 150502 97298 150554
rect 97298 150502 97350 150554
rect 97350 150502 97352 150554
rect 97296 150500 97352 150502
rect 97400 150554 97456 150556
rect 97400 150502 97402 150554
rect 97402 150502 97454 150554
rect 97454 150502 97456 150554
rect 97400 150500 97456 150502
rect 97504 150554 97560 150556
rect 97504 150502 97506 150554
rect 97506 150502 97558 150554
rect 97558 150502 97560 150554
rect 97504 150500 97560 150502
rect 128016 150554 128072 150556
rect 128016 150502 128018 150554
rect 128018 150502 128070 150554
rect 128070 150502 128072 150554
rect 128016 150500 128072 150502
rect 128120 150554 128176 150556
rect 128120 150502 128122 150554
rect 128122 150502 128174 150554
rect 128174 150502 128176 150554
rect 128120 150500 128176 150502
rect 128224 150554 128280 150556
rect 128224 150502 128226 150554
rect 128226 150502 128278 150554
rect 128278 150502 128280 150554
rect 128224 150500 128280 150502
rect 65916 149770 65972 149772
rect 65916 149718 65918 149770
rect 65918 149718 65970 149770
rect 65970 149718 65972 149770
rect 65916 149716 65972 149718
rect 66020 149770 66076 149772
rect 66020 149718 66022 149770
rect 66022 149718 66074 149770
rect 66074 149718 66076 149770
rect 66020 149716 66076 149718
rect 66124 149770 66180 149772
rect 66124 149718 66126 149770
rect 66126 149718 66178 149770
rect 66178 149718 66180 149770
rect 66124 149716 66180 149718
rect 96636 149770 96692 149772
rect 96636 149718 96638 149770
rect 96638 149718 96690 149770
rect 96690 149718 96692 149770
rect 96636 149716 96692 149718
rect 96740 149770 96796 149772
rect 96740 149718 96742 149770
rect 96742 149718 96794 149770
rect 96794 149718 96796 149770
rect 96740 149716 96796 149718
rect 96844 149770 96900 149772
rect 96844 149718 96846 149770
rect 96846 149718 96898 149770
rect 96898 149718 96900 149770
rect 96844 149716 96900 149718
rect 127356 149770 127412 149772
rect 127356 149718 127358 149770
rect 127358 149718 127410 149770
rect 127410 149718 127412 149770
rect 127356 149716 127412 149718
rect 127460 149770 127516 149772
rect 127460 149718 127462 149770
rect 127462 149718 127514 149770
rect 127514 149718 127516 149770
rect 127460 149716 127516 149718
rect 127564 149770 127620 149772
rect 127564 149718 127566 149770
rect 127566 149718 127618 149770
rect 127618 149718 127620 149770
rect 127564 149716 127620 149718
rect 158736 156826 158792 156828
rect 158736 156774 158738 156826
rect 158738 156774 158790 156826
rect 158790 156774 158792 156826
rect 158736 156772 158792 156774
rect 158840 156826 158896 156828
rect 158840 156774 158842 156826
rect 158842 156774 158894 156826
rect 158894 156774 158896 156826
rect 158840 156772 158896 156774
rect 158944 156826 159000 156828
rect 158944 156774 158946 156826
rect 158946 156774 158998 156826
rect 158998 156774 159000 156826
rect 158944 156772 159000 156774
rect 66576 148986 66632 148988
rect 66576 148934 66578 148986
rect 66578 148934 66630 148986
rect 66630 148934 66632 148986
rect 66576 148932 66632 148934
rect 66680 148986 66736 148988
rect 66680 148934 66682 148986
rect 66682 148934 66734 148986
rect 66734 148934 66736 148986
rect 66680 148932 66736 148934
rect 66784 148986 66840 148988
rect 66784 148934 66786 148986
rect 66786 148934 66838 148986
rect 66838 148934 66840 148986
rect 66784 148932 66840 148934
rect 97296 148986 97352 148988
rect 97296 148934 97298 148986
rect 97298 148934 97350 148986
rect 97350 148934 97352 148986
rect 97296 148932 97352 148934
rect 97400 148986 97456 148988
rect 97400 148934 97402 148986
rect 97402 148934 97454 148986
rect 97454 148934 97456 148986
rect 97400 148932 97456 148934
rect 97504 148986 97560 148988
rect 97504 148934 97506 148986
rect 97506 148934 97558 148986
rect 97558 148934 97560 148986
rect 97504 148932 97560 148934
rect 128016 148986 128072 148988
rect 128016 148934 128018 148986
rect 128018 148934 128070 148986
rect 128070 148934 128072 148986
rect 128016 148932 128072 148934
rect 128120 148986 128176 148988
rect 128120 148934 128122 148986
rect 128122 148934 128174 148986
rect 128174 148934 128176 148986
rect 128120 148932 128176 148934
rect 128224 148986 128280 148988
rect 128224 148934 128226 148986
rect 128226 148934 128278 148986
rect 128278 148934 128280 148986
rect 128224 148932 128280 148934
rect 65916 148202 65972 148204
rect 65916 148150 65918 148202
rect 65918 148150 65970 148202
rect 65970 148150 65972 148202
rect 65916 148148 65972 148150
rect 66020 148202 66076 148204
rect 66020 148150 66022 148202
rect 66022 148150 66074 148202
rect 66074 148150 66076 148202
rect 66020 148148 66076 148150
rect 66124 148202 66180 148204
rect 66124 148150 66126 148202
rect 66126 148150 66178 148202
rect 66178 148150 66180 148202
rect 66124 148148 66180 148150
rect 96636 148202 96692 148204
rect 96636 148150 96638 148202
rect 96638 148150 96690 148202
rect 96690 148150 96692 148202
rect 96636 148148 96692 148150
rect 96740 148202 96796 148204
rect 96740 148150 96742 148202
rect 96742 148150 96794 148202
rect 96794 148150 96796 148202
rect 96740 148148 96796 148150
rect 96844 148202 96900 148204
rect 96844 148150 96846 148202
rect 96846 148150 96898 148202
rect 96898 148150 96900 148202
rect 96844 148148 96900 148150
rect 127356 148202 127412 148204
rect 127356 148150 127358 148202
rect 127358 148150 127410 148202
rect 127410 148150 127412 148202
rect 127356 148148 127412 148150
rect 127460 148202 127516 148204
rect 127460 148150 127462 148202
rect 127462 148150 127514 148202
rect 127514 148150 127516 148202
rect 127460 148148 127516 148150
rect 127564 148202 127620 148204
rect 127564 148150 127566 148202
rect 127566 148150 127618 148202
rect 127618 148150 127620 148202
rect 127564 148148 127620 148150
rect 66576 147418 66632 147420
rect 66576 147366 66578 147418
rect 66578 147366 66630 147418
rect 66630 147366 66632 147418
rect 66576 147364 66632 147366
rect 66680 147418 66736 147420
rect 66680 147366 66682 147418
rect 66682 147366 66734 147418
rect 66734 147366 66736 147418
rect 66680 147364 66736 147366
rect 66784 147418 66840 147420
rect 66784 147366 66786 147418
rect 66786 147366 66838 147418
rect 66838 147366 66840 147418
rect 66784 147364 66840 147366
rect 97296 147418 97352 147420
rect 97296 147366 97298 147418
rect 97298 147366 97350 147418
rect 97350 147366 97352 147418
rect 97296 147364 97352 147366
rect 97400 147418 97456 147420
rect 97400 147366 97402 147418
rect 97402 147366 97454 147418
rect 97454 147366 97456 147418
rect 97400 147364 97456 147366
rect 97504 147418 97560 147420
rect 97504 147366 97506 147418
rect 97506 147366 97558 147418
rect 97558 147366 97560 147418
rect 97504 147364 97560 147366
rect 128016 147418 128072 147420
rect 128016 147366 128018 147418
rect 128018 147366 128070 147418
rect 128070 147366 128072 147418
rect 128016 147364 128072 147366
rect 128120 147418 128176 147420
rect 128120 147366 128122 147418
rect 128122 147366 128174 147418
rect 128174 147366 128176 147418
rect 128120 147364 128176 147366
rect 128224 147418 128280 147420
rect 128224 147366 128226 147418
rect 128226 147366 128278 147418
rect 128278 147366 128280 147418
rect 128224 147364 128280 147366
rect 65916 146634 65972 146636
rect 65916 146582 65918 146634
rect 65918 146582 65970 146634
rect 65970 146582 65972 146634
rect 65916 146580 65972 146582
rect 66020 146634 66076 146636
rect 66020 146582 66022 146634
rect 66022 146582 66074 146634
rect 66074 146582 66076 146634
rect 66020 146580 66076 146582
rect 66124 146634 66180 146636
rect 66124 146582 66126 146634
rect 66126 146582 66178 146634
rect 66178 146582 66180 146634
rect 66124 146580 66180 146582
rect 96636 146634 96692 146636
rect 96636 146582 96638 146634
rect 96638 146582 96690 146634
rect 96690 146582 96692 146634
rect 96636 146580 96692 146582
rect 96740 146634 96796 146636
rect 96740 146582 96742 146634
rect 96742 146582 96794 146634
rect 96794 146582 96796 146634
rect 96740 146580 96796 146582
rect 96844 146634 96900 146636
rect 96844 146582 96846 146634
rect 96846 146582 96898 146634
rect 96898 146582 96900 146634
rect 96844 146580 96900 146582
rect 127356 146634 127412 146636
rect 127356 146582 127358 146634
rect 127358 146582 127410 146634
rect 127410 146582 127412 146634
rect 127356 146580 127412 146582
rect 127460 146634 127516 146636
rect 127460 146582 127462 146634
rect 127462 146582 127514 146634
rect 127514 146582 127516 146634
rect 127460 146580 127516 146582
rect 127564 146634 127620 146636
rect 127564 146582 127566 146634
rect 127566 146582 127618 146634
rect 127618 146582 127620 146634
rect 127564 146580 127620 146582
rect 66576 145850 66632 145852
rect 66576 145798 66578 145850
rect 66578 145798 66630 145850
rect 66630 145798 66632 145850
rect 66576 145796 66632 145798
rect 66680 145850 66736 145852
rect 66680 145798 66682 145850
rect 66682 145798 66734 145850
rect 66734 145798 66736 145850
rect 66680 145796 66736 145798
rect 66784 145850 66840 145852
rect 66784 145798 66786 145850
rect 66786 145798 66838 145850
rect 66838 145798 66840 145850
rect 66784 145796 66840 145798
rect 97296 145850 97352 145852
rect 97296 145798 97298 145850
rect 97298 145798 97350 145850
rect 97350 145798 97352 145850
rect 97296 145796 97352 145798
rect 97400 145850 97456 145852
rect 97400 145798 97402 145850
rect 97402 145798 97454 145850
rect 97454 145798 97456 145850
rect 97400 145796 97456 145798
rect 97504 145850 97560 145852
rect 97504 145798 97506 145850
rect 97506 145798 97558 145850
rect 97558 145798 97560 145850
rect 97504 145796 97560 145798
rect 128016 145850 128072 145852
rect 128016 145798 128018 145850
rect 128018 145798 128070 145850
rect 128070 145798 128072 145850
rect 128016 145796 128072 145798
rect 128120 145850 128176 145852
rect 128120 145798 128122 145850
rect 128122 145798 128174 145850
rect 128174 145798 128176 145850
rect 128120 145796 128176 145798
rect 128224 145850 128280 145852
rect 128224 145798 128226 145850
rect 128226 145798 128278 145850
rect 128278 145798 128280 145850
rect 128224 145796 128280 145798
rect 65916 145066 65972 145068
rect 65916 145014 65918 145066
rect 65918 145014 65970 145066
rect 65970 145014 65972 145066
rect 65916 145012 65972 145014
rect 66020 145066 66076 145068
rect 66020 145014 66022 145066
rect 66022 145014 66074 145066
rect 66074 145014 66076 145066
rect 66020 145012 66076 145014
rect 66124 145066 66180 145068
rect 66124 145014 66126 145066
rect 66126 145014 66178 145066
rect 66178 145014 66180 145066
rect 66124 145012 66180 145014
rect 96636 145066 96692 145068
rect 96636 145014 96638 145066
rect 96638 145014 96690 145066
rect 96690 145014 96692 145066
rect 96636 145012 96692 145014
rect 96740 145066 96796 145068
rect 96740 145014 96742 145066
rect 96742 145014 96794 145066
rect 96794 145014 96796 145066
rect 96740 145012 96796 145014
rect 96844 145066 96900 145068
rect 96844 145014 96846 145066
rect 96846 145014 96898 145066
rect 96898 145014 96900 145066
rect 96844 145012 96900 145014
rect 127356 145066 127412 145068
rect 127356 145014 127358 145066
rect 127358 145014 127410 145066
rect 127410 145014 127412 145066
rect 127356 145012 127412 145014
rect 127460 145066 127516 145068
rect 127460 145014 127462 145066
rect 127462 145014 127514 145066
rect 127514 145014 127516 145066
rect 127460 145012 127516 145014
rect 127564 145066 127620 145068
rect 127564 145014 127566 145066
rect 127566 145014 127618 145066
rect 127618 145014 127620 145066
rect 127564 145012 127620 145014
rect 132972 46956 133028 47012
rect 158076 156042 158132 156044
rect 158076 155990 158078 156042
rect 158078 155990 158130 156042
rect 158130 155990 158132 156042
rect 158076 155988 158132 155990
rect 158180 156042 158236 156044
rect 158180 155990 158182 156042
rect 158182 155990 158234 156042
rect 158234 155990 158236 156042
rect 158180 155988 158236 155990
rect 158284 156042 158340 156044
rect 158284 155990 158286 156042
rect 158286 155990 158338 156042
rect 158338 155990 158340 156042
rect 158284 155988 158340 155990
rect 189456 156826 189512 156828
rect 189456 156774 189458 156826
rect 189458 156774 189510 156826
rect 189510 156774 189512 156826
rect 189456 156772 189512 156774
rect 189560 156826 189616 156828
rect 189560 156774 189562 156826
rect 189562 156774 189614 156826
rect 189614 156774 189616 156826
rect 189560 156772 189616 156774
rect 189664 156826 189720 156828
rect 189664 156774 189666 156826
rect 189666 156774 189718 156826
rect 189718 156774 189720 156826
rect 189664 156772 189720 156774
rect 188796 156042 188852 156044
rect 188796 155990 188798 156042
rect 188798 155990 188850 156042
rect 188850 155990 188852 156042
rect 188796 155988 188852 155990
rect 188900 156042 188956 156044
rect 188900 155990 188902 156042
rect 188902 155990 188954 156042
rect 188954 155990 188956 156042
rect 188900 155988 188956 155990
rect 189004 156042 189060 156044
rect 189004 155990 189006 156042
rect 189006 155990 189058 156042
rect 189058 155990 189060 156042
rect 189004 155988 189060 155990
rect 194236 155820 194292 155876
rect 194908 155820 194964 155876
rect 158736 155258 158792 155260
rect 158736 155206 158738 155258
rect 158738 155206 158790 155258
rect 158790 155206 158792 155258
rect 158736 155204 158792 155206
rect 158840 155258 158896 155260
rect 158840 155206 158842 155258
rect 158842 155206 158894 155258
rect 158894 155206 158896 155258
rect 158840 155204 158896 155206
rect 158944 155258 159000 155260
rect 158944 155206 158946 155258
rect 158946 155206 158998 155258
rect 158998 155206 159000 155258
rect 158944 155204 159000 155206
rect 158076 154474 158132 154476
rect 158076 154422 158078 154474
rect 158078 154422 158130 154474
rect 158130 154422 158132 154474
rect 158076 154420 158132 154422
rect 158180 154474 158236 154476
rect 158180 154422 158182 154474
rect 158182 154422 158234 154474
rect 158234 154422 158236 154474
rect 158180 154420 158236 154422
rect 158284 154474 158340 154476
rect 158284 154422 158286 154474
rect 158286 154422 158338 154474
rect 158338 154422 158340 154474
rect 158284 154420 158340 154422
rect 158736 153690 158792 153692
rect 158736 153638 158738 153690
rect 158738 153638 158790 153690
rect 158790 153638 158792 153690
rect 158736 153636 158792 153638
rect 158840 153690 158896 153692
rect 158840 153638 158842 153690
rect 158842 153638 158894 153690
rect 158894 153638 158896 153690
rect 158840 153636 158896 153638
rect 158944 153690 159000 153692
rect 158944 153638 158946 153690
rect 158946 153638 158998 153690
rect 158998 153638 159000 153690
rect 158944 153636 159000 153638
rect 158076 152906 158132 152908
rect 158076 152854 158078 152906
rect 158078 152854 158130 152906
rect 158130 152854 158132 152906
rect 158076 152852 158132 152854
rect 158180 152906 158236 152908
rect 158180 152854 158182 152906
rect 158182 152854 158234 152906
rect 158234 152854 158236 152906
rect 158180 152852 158236 152854
rect 158284 152906 158340 152908
rect 158284 152854 158286 152906
rect 158286 152854 158338 152906
rect 158338 152854 158340 152906
rect 158284 152852 158340 152854
rect 158736 152122 158792 152124
rect 158736 152070 158738 152122
rect 158738 152070 158790 152122
rect 158790 152070 158792 152122
rect 158736 152068 158792 152070
rect 158840 152122 158896 152124
rect 158840 152070 158842 152122
rect 158842 152070 158894 152122
rect 158894 152070 158896 152122
rect 158840 152068 158896 152070
rect 158944 152122 159000 152124
rect 158944 152070 158946 152122
rect 158946 152070 158998 152122
rect 158998 152070 159000 152122
rect 158944 152068 159000 152070
rect 158076 151338 158132 151340
rect 158076 151286 158078 151338
rect 158078 151286 158130 151338
rect 158130 151286 158132 151338
rect 158076 151284 158132 151286
rect 158180 151338 158236 151340
rect 158180 151286 158182 151338
rect 158182 151286 158234 151338
rect 158234 151286 158236 151338
rect 158180 151284 158236 151286
rect 158284 151338 158340 151340
rect 158284 151286 158286 151338
rect 158286 151286 158338 151338
rect 158338 151286 158340 151338
rect 158284 151284 158340 151286
rect 158736 150554 158792 150556
rect 158736 150502 158738 150554
rect 158738 150502 158790 150554
rect 158790 150502 158792 150554
rect 158736 150500 158792 150502
rect 158840 150554 158896 150556
rect 158840 150502 158842 150554
rect 158842 150502 158894 150554
rect 158894 150502 158896 150554
rect 158840 150500 158896 150502
rect 158944 150554 159000 150556
rect 158944 150502 158946 150554
rect 158946 150502 158998 150554
rect 158998 150502 159000 150554
rect 158944 150500 159000 150502
rect 158076 149770 158132 149772
rect 158076 149718 158078 149770
rect 158078 149718 158130 149770
rect 158130 149718 158132 149770
rect 158076 149716 158132 149718
rect 158180 149770 158236 149772
rect 158180 149718 158182 149770
rect 158182 149718 158234 149770
rect 158234 149718 158236 149770
rect 158180 149716 158236 149718
rect 158284 149770 158340 149772
rect 158284 149718 158286 149770
rect 158286 149718 158338 149770
rect 158338 149718 158340 149770
rect 158284 149716 158340 149718
rect 189456 155258 189512 155260
rect 189456 155206 189458 155258
rect 189458 155206 189510 155258
rect 189510 155206 189512 155258
rect 189456 155204 189512 155206
rect 189560 155258 189616 155260
rect 189560 155206 189562 155258
rect 189562 155206 189614 155258
rect 189614 155206 189616 155258
rect 189560 155204 189616 155206
rect 189664 155258 189720 155260
rect 189664 155206 189666 155258
rect 189666 155206 189718 155258
rect 189718 155206 189720 155258
rect 189664 155204 189720 155206
rect 188796 154474 188852 154476
rect 188796 154422 188798 154474
rect 188798 154422 188850 154474
rect 188850 154422 188852 154474
rect 188796 154420 188852 154422
rect 188900 154474 188956 154476
rect 188900 154422 188902 154474
rect 188902 154422 188954 154474
rect 188954 154422 188956 154474
rect 188900 154420 188956 154422
rect 189004 154474 189060 154476
rect 189004 154422 189006 154474
rect 189006 154422 189058 154474
rect 189058 154422 189060 154474
rect 189004 154420 189060 154422
rect 189456 153690 189512 153692
rect 189456 153638 189458 153690
rect 189458 153638 189510 153690
rect 189510 153638 189512 153690
rect 189456 153636 189512 153638
rect 189560 153690 189616 153692
rect 189560 153638 189562 153690
rect 189562 153638 189614 153690
rect 189614 153638 189616 153690
rect 189560 153636 189616 153638
rect 189664 153690 189720 153692
rect 189664 153638 189666 153690
rect 189666 153638 189718 153690
rect 189718 153638 189720 153690
rect 189664 153636 189720 153638
rect 188796 152906 188852 152908
rect 188796 152854 188798 152906
rect 188798 152854 188850 152906
rect 188850 152854 188852 152906
rect 188796 152852 188852 152854
rect 188900 152906 188956 152908
rect 188900 152854 188902 152906
rect 188902 152854 188954 152906
rect 188954 152854 188956 152906
rect 188900 152852 188956 152854
rect 189004 152906 189060 152908
rect 189004 152854 189006 152906
rect 189006 152854 189058 152906
rect 189058 152854 189060 152906
rect 189004 152852 189060 152854
rect 189456 152122 189512 152124
rect 189456 152070 189458 152122
rect 189458 152070 189510 152122
rect 189510 152070 189512 152122
rect 189456 152068 189512 152070
rect 189560 152122 189616 152124
rect 189560 152070 189562 152122
rect 189562 152070 189614 152122
rect 189614 152070 189616 152122
rect 189560 152068 189616 152070
rect 189664 152122 189720 152124
rect 189664 152070 189666 152122
rect 189666 152070 189718 152122
rect 189718 152070 189720 152122
rect 189664 152068 189720 152070
rect 188796 151338 188852 151340
rect 188796 151286 188798 151338
rect 188798 151286 188850 151338
rect 188850 151286 188852 151338
rect 188796 151284 188852 151286
rect 188900 151338 188956 151340
rect 188900 151286 188902 151338
rect 188902 151286 188954 151338
rect 188954 151286 188956 151338
rect 188900 151284 188956 151286
rect 189004 151338 189060 151340
rect 189004 151286 189006 151338
rect 189006 151286 189058 151338
rect 189058 151286 189060 151338
rect 189004 151284 189060 151286
rect 189456 150554 189512 150556
rect 189456 150502 189458 150554
rect 189458 150502 189510 150554
rect 189510 150502 189512 150554
rect 189456 150500 189512 150502
rect 189560 150554 189616 150556
rect 189560 150502 189562 150554
rect 189562 150502 189614 150554
rect 189614 150502 189616 150554
rect 189560 150500 189616 150502
rect 189664 150554 189720 150556
rect 189664 150502 189666 150554
rect 189666 150502 189718 150554
rect 189718 150502 189720 150554
rect 189664 150500 189720 150502
rect 188796 149770 188852 149772
rect 188796 149718 188798 149770
rect 188798 149718 188850 149770
rect 188850 149718 188852 149770
rect 188796 149716 188852 149718
rect 188900 149770 188956 149772
rect 188900 149718 188902 149770
rect 188902 149718 188954 149770
rect 188954 149718 188956 149770
rect 188900 149716 188956 149718
rect 189004 149770 189060 149772
rect 189004 149718 189006 149770
rect 189006 149718 189058 149770
rect 189058 149718 189060 149770
rect 189004 149716 189060 149718
rect 158736 148986 158792 148988
rect 158736 148934 158738 148986
rect 158738 148934 158790 148986
rect 158790 148934 158792 148986
rect 158736 148932 158792 148934
rect 158840 148986 158896 148988
rect 158840 148934 158842 148986
rect 158842 148934 158894 148986
rect 158894 148934 158896 148986
rect 158840 148932 158896 148934
rect 158944 148986 159000 148988
rect 158944 148934 158946 148986
rect 158946 148934 158998 148986
rect 158998 148934 159000 148986
rect 158944 148932 159000 148934
rect 158076 148202 158132 148204
rect 158076 148150 158078 148202
rect 158078 148150 158130 148202
rect 158130 148150 158132 148202
rect 158076 148148 158132 148150
rect 158180 148202 158236 148204
rect 158180 148150 158182 148202
rect 158182 148150 158234 148202
rect 158234 148150 158236 148202
rect 158180 148148 158236 148150
rect 158284 148202 158340 148204
rect 158284 148150 158286 148202
rect 158286 148150 158338 148202
rect 158338 148150 158340 148202
rect 158284 148148 158340 148150
rect 158736 147418 158792 147420
rect 158736 147366 158738 147418
rect 158738 147366 158790 147418
rect 158790 147366 158792 147418
rect 158736 147364 158792 147366
rect 158840 147418 158896 147420
rect 158840 147366 158842 147418
rect 158842 147366 158894 147418
rect 158894 147366 158896 147418
rect 158840 147364 158896 147366
rect 158944 147418 159000 147420
rect 158944 147366 158946 147418
rect 158946 147366 158998 147418
rect 158998 147366 159000 147418
rect 158944 147364 159000 147366
rect 158076 146634 158132 146636
rect 158076 146582 158078 146634
rect 158078 146582 158130 146634
rect 158130 146582 158132 146634
rect 158076 146580 158132 146582
rect 158180 146634 158236 146636
rect 158180 146582 158182 146634
rect 158182 146582 158234 146634
rect 158234 146582 158236 146634
rect 158180 146580 158236 146582
rect 158284 146634 158340 146636
rect 158284 146582 158286 146634
rect 158286 146582 158338 146634
rect 158338 146582 158340 146634
rect 158284 146580 158340 146582
rect 158736 145850 158792 145852
rect 158736 145798 158738 145850
rect 158738 145798 158790 145850
rect 158790 145798 158792 145850
rect 158736 145796 158792 145798
rect 158840 145850 158896 145852
rect 158840 145798 158842 145850
rect 158842 145798 158894 145850
rect 158894 145798 158896 145850
rect 158840 145796 158896 145798
rect 158944 145850 159000 145852
rect 158944 145798 158946 145850
rect 158946 145798 158998 145850
rect 158998 145798 159000 145850
rect 158944 145796 159000 145798
rect 158076 145066 158132 145068
rect 158076 145014 158078 145066
rect 158078 145014 158130 145066
rect 158130 145014 158132 145066
rect 158076 145012 158132 145014
rect 158180 145066 158236 145068
rect 158180 145014 158182 145066
rect 158182 145014 158234 145066
rect 158234 145014 158236 145066
rect 158180 145012 158236 145014
rect 158284 145066 158340 145068
rect 158284 145014 158286 145066
rect 158286 145014 158338 145066
rect 158338 145014 158340 145066
rect 158284 145012 158340 145014
rect 156380 46956 156436 47012
rect 132972 45724 133028 45780
rect 71932 41244 71988 41300
rect 67676 41020 67732 41076
rect 65100 22316 65156 22372
rect 59052 19852 59108 19908
rect 75516 41132 75572 41188
rect 71932 22316 71988 22372
rect 67676 21756 67732 21812
rect 68796 21756 68852 21812
rect 67788 20412 67844 20468
rect 66576 17274 66632 17276
rect 66576 17222 66578 17274
rect 66578 17222 66630 17274
rect 66630 17222 66632 17274
rect 66576 17220 66632 17222
rect 66680 17274 66736 17276
rect 66680 17222 66682 17274
rect 66682 17222 66734 17274
rect 66734 17222 66736 17274
rect 66680 17220 66736 17222
rect 66784 17274 66840 17276
rect 66784 17222 66786 17274
rect 66786 17222 66838 17274
rect 66838 17222 66840 17274
rect 66784 17220 66840 17222
rect 85148 40908 85204 40964
rect 132972 38108 133028 38164
rect 156380 45724 156436 45780
rect 189456 148986 189512 148988
rect 189456 148934 189458 148986
rect 189458 148934 189510 148986
rect 189510 148934 189512 148986
rect 189456 148932 189512 148934
rect 189560 148986 189616 148988
rect 189560 148934 189562 148986
rect 189562 148934 189614 148986
rect 189614 148934 189616 148986
rect 189560 148932 189616 148934
rect 189664 148986 189720 148988
rect 189664 148934 189666 148986
rect 189666 148934 189718 148986
rect 189718 148934 189720 148986
rect 189664 148932 189720 148934
rect 188796 148202 188852 148204
rect 188796 148150 188798 148202
rect 188798 148150 188850 148202
rect 188850 148150 188852 148202
rect 188796 148148 188852 148150
rect 188900 148202 188956 148204
rect 188900 148150 188902 148202
rect 188902 148150 188954 148202
rect 188954 148150 188956 148202
rect 188900 148148 188956 148150
rect 189004 148202 189060 148204
rect 189004 148150 189006 148202
rect 189006 148150 189058 148202
rect 189058 148150 189060 148202
rect 189004 148148 189060 148150
rect 189456 147418 189512 147420
rect 189456 147366 189458 147418
rect 189458 147366 189510 147418
rect 189510 147366 189512 147418
rect 189456 147364 189512 147366
rect 189560 147418 189616 147420
rect 189560 147366 189562 147418
rect 189562 147366 189614 147418
rect 189614 147366 189616 147418
rect 189560 147364 189616 147366
rect 189664 147418 189720 147420
rect 189664 147366 189666 147418
rect 189666 147366 189718 147418
rect 189718 147366 189720 147418
rect 189664 147364 189720 147366
rect 188796 146634 188852 146636
rect 188796 146582 188798 146634
rect 188798 146582 188850 146634
rect 188850 146582 188852 146634
rect 188796 146580 188852 146582
rect 188900 146634 188956 146636
rect 188900 146582 188902 146634
rect 188902 146582 188954 146634
rect 188954 146582 188956 146634
rect 188900 146580 188956 146582
rect 189004 146634 189060 146636
rect 189004 146582 189006 146634
rect 189006 146582 189058 146634
rect 189058 146582 189060 146634
rect 189004 146580 189060 146582
rect 189456 145850 189512 145852
rect 189456 145798 189458 145850
rect 189458 145798 189510 145850
rect 189510 145798 189512 145850
rect 189456 145796 189512 145798
rect 189560 145850 189616 145852
rect 189560 145798 189562 145850
rect 189562 145798 189614 145850
rect 189614 145798 189616 145850
rect 189560 145796 189616 145798
rect 189664 145850 189720 145852
rect 189664 145798 189666 145850
rect 189666 145798 189718 145850
rect 189718 145798 189720 145850
rect 189664 145796 189720 145798
rect 188796 145066 188852 145068
rect 188796 145014 188798 145066
rect 188798 145014 188850 145066
rect 188850 145014 188852 145066
rect 188796 145012 188852 145014
rect 188900 145066 188956 145068
rect 188900 145014 188902 145066
rect 188902 145014 188954 145066
rect 188954 145014 188956 145066
rect 188900 145012 188956 145014
rect 189004 145066 189060 145068
rect 189004 145014 189006 145066
rect 189006 145014 189058 145066
rect 189058 145014 189060 145066
rect 189004 145012 189060 145014
rect 189456 144282 189512 144284
rect 189456 144230 189458 144282
rect 189458 144230 189510 144282
rect 189510 144230 189512 144282
rect 189456 144228 189512 144230
rect 189560 144282 189616 144284
rect 189560 144230 189562 144282
rect 189562 144230 189614 144282
rect 189614 144230 189616 144282
rect 189560 144228 189616 144230
rect 189664 144282 189720 144284
rect 189664 144230 189666 144282
rect 189666 144230 189718 144282
rect 189718 144230 189720 144282
rect 189664 144228 189720 144230
rect 188796 143498 188852 143500
rect 188796 143446 188798 143498
rect 188798 143446 188850 143498
rect 188850 143446 188852 143498
rect 188796 143444 188852 143446
rect 188900 143498 188956 143500
rect 188900 143446 188902 143498
rect 188902 143446 188954 143498
rect 188954 143446 188956 143498
rect 188900 143444 188956 143446
rect 189004 143498 189060 143500
rect 189004 143446 189006 143498
rect 189006 143446 189058 143498
rect 189058 143446 189060 143498
rect 189004 143444 189060 143446
rect 189456 142714 189512 142716
rect 189456 142662 189458 142714
rect 189458 142662 189510 142714
rect 189510 142662 189512 142714
rect 189456 142660 189512 142662
rect 189560 142714 189616 142716
rect 189560 142662 189562 142714
rect 189562 142662 189614 142714
rect 189614 142662 189616 142714
rect 189560 142660 189616 142662
rect 189664 142714 189720 142716
rect 189664 142662 189666 142714
rect 189666 142662 189718 142714
rect 189718 142662 189720 142714
rect 189664 142660 189720 142662
rect 188796 141930 188852 141932
rect 188796 141878 188798 141930
rect 188798 141878 188850 141930
rect 188850 141878 188852 141930
rect 188796 141876 188852 141878
rect 188900 141930 188956 141932
rect 188900 141878 188902 141930
rect 188902 141878 188954 141930
rect 188954 141878 188956 141930
rect 188900 141876 188956 141878
rect 189004 141930 189060 141932
rect 189004 141878 189006 141930
rect 189006 141878 189058 141930
rect 189058 141878 189060 141930
rect 189004 141876 189060 141878
rect 189456 141146 189512 141148
rect 189456 141094 189458 141146
rect 189458 141094 189510 141146
rect 189510 141094 189512 141146
rect 189456 141092 189512 141094
rect 189560 141146 189616 141148
rect 189560 141094 189562 141146
rect 189562 141094 189614 141146
rect 189614 141094 189616 141146
rect 189560 141092 189616 141094
rect 189664 141146 189720 141148
rect 189664 141094 189666 141146
rect 189666 141094 189718 141146
rect 189718 141094 189720 141146
rect 189664 141092 189720 141094
rect 188796 140362 188852 140364
rect 188796 140310 188798 140362
rect 188798 140310 188850 140362
rect 188850 140310 188852 140362
rect 188796 140308 188852 140310
rect 188900 140362 188956 140364
rect 188900 140310 188902 140362
rect 188902 140310 188954 140362
rect 188954 140310 188956 140362
rect 188900 140308 188956 140310
rect 189004 140362 189060 140364
rect 189004 140310 189006 140362
rect 189006 140310 189058 140362
rect 189058 140310 189060 140362
rect 189004 140308 189060 140310
rect 189456 139578 189512 139580
rect 189456 139526 189458 139578
rect 189458 139526 189510 139578
rect 189510 139526 189512 139578
rect 189456 139524 189512 139526
rect 189560 139578 189616 139580
rect 189560 139526 189562 139578
rect 189562 139526 189614 139578
rect 189614 139526 189616 139578
rect 189560 139524 189616 139526
rect 189664 139578 189720 139580
rect 189664 139526 189666 139578
rect 189666 139526 189718 139578
rect 189718 139526 189720 139578
rect 189664 139524 189720 139526
rect 188796 138794 188852 138796
rect 188796 138742 188798 138794
rect 188798 138742 188850 138794
rect 188850 138742 188852 138794
rect 188796 138740 188852 138742
rect 188900 138794 188956 138796
rect 188900 138742 188902 138794
rect 188902 138742 188954 138794
rect 188954 138742 188956 138794
rect 188900 138740 188956 138742
rect 189004 138794 189060 138796
rect 189004 138742 189006 138794
rect 189006 138742 189058 138794
rect 189058 138742 189060 138794
rect 189004 138740 189060 138742
rect 189456 138010 189512 138012
rect 189456 137958 189458 138010
rect 189458 137958 189510 138010
rect 189510 137958 189512 138010
rect 189456 137956 189512 137958
rect 189560 138010 189616 138012
rect 189560 137958 189562 138010
rect 189562 137958 189614 138010
rect 189614 137958 189616 138010
rect 189560 137956 189616 137958
rect 189664 138010 189720 138012
rect 189664 137958 189666 138010
rect 189666 137958 189718 138010
rect 189718 137958 189720 138010
rect 189664 137956 189720 137958
rect 188796 137226 188852 137228
rect 188796 137174 188798 137226
rect 188798 137174 188850 137226
rect 188850 137174 188852 137226
rect 188796 137172 188852 137174
rect 188900 137226 188956 137228
rect 188900 137174 188902 137226
rect 188902 137174 188954 137226
rect 188954 137174 188956 137226
rect 188900 137172 188956 137174
rect 189004 137226 189060 137228
rect 189004 137174 189006 137226
rect 189006 137174 189058 137226
rect 189058 137174 189060 137226
rect 189004 137172 189060 137174
rect 189456 136442 189512 136444
rect 189456 136390 189458 136442
rect 189458 136390 189510 136442
rect 189510 136390 189512 136442
rect 189456 136388 189512 136390
rect 189560 136442 189616 136444
rect 189560 136390 189562 136442
rect 189562 136390 189614 136442
rect 189614 136390 189616 136442
rect 189560 136388 189616 136390
rect 189664 136442 189720 136444
rect 189664 136390 189666 136442
rect 189666 136390 189718 136442
rect 189718 136390 189720 136442
rect 189664 136388 189720 136390
rect 188796 135658 188852 135660
rect 188796 135606 188798 135658
rect 188798 135606 188850 135658
rect 188850 135606 188852 135658
rect 188796 135604 188852 135606
rect 188900 135658 188956 135660
rect 188900 135606 188902 135658
rect 188902 135606 188954 135658
rect 188954 135606 188956 135658
rect 188900 135604 188956 135606
rect 189004 135658 189060 135660
rect 189004 135606 189006 135658
rect 189006 135606 189058 135658
rect 189058 135606 189060 135658
rect 189004 135604 189060 135606
rect 189456 134874 189512 134876
rect 189456 134822 189458 134874
rect 189458 134822 189510 134874
rect 189510 134822 189512 134874
rect 189456 134820 189512 134822
rect 189560 134874 189616 134876
rect 189560 134822 189562 134874
rect 189562 134822 189614 134874
rect 189614 134822 189616 134874
rect 189560 134820 189616 134822
rect 189664 134874 189720 134876
rect 189664 134822 189666 134874
rect 189666 134822 189718 134874
rect 189718 134822 189720 134874
rect 189664 134820 189720 134822
rect 188796 134090 188852 134092
rect 188796 134038 188798 134090
rect 188798 134038 188850 134090
rect 188850 134038 188852 134090
rect 188796 134036 188852 134038
rect 188900 134090 188956 134092
rect 188900 134038 188902 134090
rect 188902 134038 188954 134090
rect 188954 134038 188956 134090
rect 188900 134036 188956 134038
rect 189004 134090 189060 134092
rect 189004 134038 189006 134090
rect 189006 134038 189058 134090
rect 189058 134038 189060 134090
rect 189004 134036 189060 134038
rect 189456 133306 189512 133308
rect 189456 133254 189458 133306
rect 189458 133254 189510 133306
rect 189510 133254 189512 133306
rect 189456 133252 189512 133254
rect 189560 133306 189616 133308
rect 189560 133254 189562 133306
rect 189562 133254 189614 133306
rect 189614 133254 189616 133306
rect 189560 133252 189616 133254
rect 189664 133306 189720 133308
rect 189664 133254 189666 133306
rect 189666 133254 189718 133306
rect 189718 133254 189720 133306
rect 189664 133252 189720 133254
rect 188796 132522 188852 132524
rect 188796 132470 188798 132522
rect 188798 132470 188850 132522
rect 188850 132470 188852 132522
rect 188796 132468 188852 132470
rect 188900 132522 188956 132524
rect 188900 132470 188902 132522
rect 188902 132470 188954 132522
rect 188954 132470 188956 132522
rect 188900 132468 188956 132470
rect 189004 132522 189060 132524
rect 189004 132470 189006 132522
rect 189006 132470 189058 132522
rect 189058 132470 189060 132522
rect 189004 132468 189060 132470
rect 189456 131738 189512 131740
rect 189456 131686 189458 131738
rect 189458 131686 189510 131738
rect 189510 131686 189512 131738
rect 189456 131684 189512 131686
rect 189560 131738 189616 131740
rect 189560 131686 189562 131738
rect 189562 131686 189614 131738
rect 189614 131686 189616 131738
rect 189560 131684 189616 131686
rect 189664 131738 189720 131740
rect 189664 131686 189666 131738
rect 189666 131686 189718 131738
rect 189718 131686 189720 131738
rect 189664 131684 189720 131686
rect 188796 130954 188852 130956
rect 188796 130902 188798 130954
rect 188798 130902 188850 130954
rect 188850 130902 188852 130954
rect 188796 130900 188852 130902
rect 188900 130954 188956 130956
rect 188900 130902 188902 130954
rect 188902 130902 188954 130954
rect 188954 130902 188956 130954
rect 188900 130900 188956 130902
rect 189004 130954 189060 130956
rect 189004 130902 189006 130954
rect 189006 130902 189058 130954
rect 189058 130902 189060 130954
rect 189004 130900 189060 130902
rect 189456 130170 189512 130172
rect 189456 130118 189458 130170
rect 189458 130118 189510 130170
rect 189510 130118 189512 130170
rect 189456 130116 189512 130118
rect 189560 130170 189616 130172
rect 189560 130118 189562 130170
rect 189562 130118 189614 130170
rect 189614 130118 189616 130170
rect 189560 130116 189616 130118
rect 189664 130170 189720 130172
rect 189664 130118 189666 130170
rect 189666 130118 189718 130170
rect 189718 130118 189720 130170
rect 189664 130116 189720 130118
rect 188796 129386 188852 129388
rect 188796 129334 188798 129386
rect 188798 129334 188850 129386
rect 188850 129334 188852 129386
rect 188796 129332 188852 129334
rect 188900 129386 188956 129388
rect 188900 129334 188902 129386
rect 188902 129334 188954 129386
rect 188954 129334 188956 129386
rect 188900 129332 188956 129334
rect 189004 129386 189060 129388
rect 189004 129334 189006 129386
rect 189006 129334 189058 129386
rect 189058 129334 189060 129386
rect 189004 129332 189060 129334
rect 189456 128602 189512 128604
rect 189456 128550 189458 128602
rect 189458 128550 189510 128602
rect 189510 128550 189512 128602
rect 189456 128548 189512 128550
rect 189560 128602 189616 128604
rect 189560 128550 189562 128602
rect 189562 128550 189614 128602
rect 189614 128550 189616 128602
rect 189560 128548 189616 128550
rect 189664 128602 189720 128604
rect 189664 128550 189666 128602
rect 189666 128550 189718 128602
rect 189718 128550 189720 128602
rect 189664 128548 189720 128550
rect 188796 127818 188852 127820
rect 188796 127766 188798 127818
rect 188798 127766 188850 127818
rect 188850 127766 188852 127818
rect 188796 127764 188852 127766
rect 188900 127818 188956 127820
rect 188900 127766 188902 127818
rect 188902 127766 188954 127818
rect 188954 127766 188956 127818
rect 188900 127764 188956 127766
rect 189004 127818 189060 127820
rect 189004 127766 189006 127818
rect 189006 127766 189058 127818
rect 189058 127766 189060 127818
rect 189004 127764 189060 127766
rect 189456 127034 189512 127036
rect 189456 126982 189458 127034
rect 189458 126982 189510 127034
rect 189510 126982 189512 127034
rect 189456 126980 189512 126982
rect 189560 127034 189616 127036
rect 189560 126982 189562 127034
rect 189562 126982 189614 127034
rect 189614 126982 189616 127034
rect 189560 126980 189616 126982
rect 189664 127034 189720 127036
rect 189664 126982 189666 127034
rect 189666 126982 189718 127034
rect 189718 126982 189720 127034
rect 189664 126980 189720 126982
rect 188796 126250 188852 126252
rect 188796 126198 188798 126250
rect 188798 126198 188850 126250
rect 188850 126198 188852 126250
rect 188796 126196 188852 126198
rect 188900 126250 188956 126252
rect 188900 126198 188902 126250
rect 188902 126198 188954 126250
rect 188954 126198 188956 126250
rect 188900 126196 188956 126198
rect 189004 126250 189060 126252
rect 189004 126198 189006 126250
rect 189006 126198 189058 126250
rect 189058 126198 189060 126250
rect 189004 126196 189060 126198
rect 189456 125466 189512 125468
rect 189456 125414 189458 125466
rect 189458 125414 189510 125466
rect 189510 125414 189512 125466
rect 189456 125412 189512 125414
rect 189560 125466 189616 125468
rect 189560 125414 189562 125466
rect 189562 125414 189614 125466
rect 189614 125414 189616 125466
rect 189560 125412 189616 125414
rect 189664 125466 189720 125468
rect 189664 125414 189666 125466
rect 189666 125414 189718 125466
rect 189718 125414 189720 125466
rect 189664 125412 189720 125414
rect 188796 124682 188852 124684
rect 188796 124630 188798 124682
rect 188798 124630 188850 124682
rect 188850 124630 188852 124682
rect 188796 124628 188852 124630
rect 188900 124682 188956 124684
rect 188900 124630 188902 124682
rect 188902 124630 188954 124682
rect 188954 124630 188956 124682
rect 188900 124628 188956 124630
rect 189004 124682 189060 124684
rect 189004 124630 189006 124682
rect 189006 124630 189058 124682
rect 189058 124630 189060 124682
rect 189004 124628 189060 124630
rect 189456 123898 189512 123900
rect 189456 123846 189458 123898
rect 189458 123846 189510 123898
rect 189510 123846 189512 123898
rect 189456 123844 189512 123846
rect 189560 123898 189616 123900
rect 189560 123846 189562 123898
rect 189562 123846 189614 123898
rect 189614 123846 189616 123898
rect 189560 123844 189616 123846
rect 189664 123898 189720 123900
rect 189664 123846 189666 123898
rect 189666 123846 189718 123898
rect 189718 123846 189720 123898
rect 189664 123844 189720 123846
rect 188796 123114 188852 123116
rect 188796 123062 188798 123114
rect 188798 123062 188850 123114
rect 188850 123062 188852 123114
rect 188796 123060 188852 123062
rect 188900 123114 188956 123116
rect 188900 123062 188902 123114
rect 188902 123062 188954 123114
rect 188954 123062 188956 123114
rect 188900 123060 188956 123062
rect 189004 123114 189060 123116
rect 189004 123062 189006 123114
rect 189006 123062 189058 123114
rect 189058 123062 189060 123114
rect 189004 123060 189060 123062
rect 189456 122330 189512 122332
rect 189456 122278 189458 122330
rect 189458 122278 189510 122330
rect 189510 122278 189512 122330
rect 189456 122276 189512 122278
rect 189560 122330 189616 122332
rect 189560 122278 189562 122330
rect 189562 122278 189614 122330
rect 189614 122278 189616 122330
rect 189560 122276 189616 122278
rect 189664 122330 189720 122332
rect 189664 122278 189666 122330
rect 189666 122278 189718 122330
rect 189718 122278 189720 122330
rect 189664 122276 189720 122278
rect 188796 121546 188852 121548
rect 188796 121494 188798 121546
rect 188798 121494 188850 121546
rect 188850 121494 188852 121546
rect 188796 121492 188852 121494
rect 188900 121546 188956 121548
rect 188900 121494 188902 121546
rect 188902 121494 188954 121546
rect 188954 121494 188956 121546
rect 188900 121492 188956 121494
rect 189004 121546 189060 121548
rect 189004 121494 189006 121546
rect 189006 121494 189058 121546
rect 189058 121494 189060 121546
rect 189004 121492 189060 121494
rect 189456 120762 189512 120764
rect 189456 120710 189458 120762
rect 189458 120710 189510 120762
rect 189510 120710 189512 120762
rect 189456 120708 189512 120710
rect 189560 120762 189616 120764
rect 189560 120710 189562 120762
rect 189562 120710 189614 120762
rect 189614 120710 189616 120762
rect 189560 120708 189616 120710
rect 189664 120762 189720 120764
rect 189664 120710 189666 120762
rect 189666 120710 189718 120762
rect 189718 120710 189720 120762
rect 189664 120708 189720 120710
rect 188796 119978 188852 119980
rect 188796 119926 188798 119978
rect 188798 119926 188850 119978
rect 188850 119926 188852 119978
rect 188796 119924 188852 119926
rect 188900 119978 188956 119980
rect 188900 119926 188902 119978
rect 188902 119926 188954 119978
rect 188954 119926 188956 119978
rect 188900 119924 188956 119926
rect 189004 119978 189060 119980
rect 189004 119926 189006 119978
rect 189006 119926 189058 119978
rect 189058 119926 189060 119978
rect 189004 119924 189060 119926
rect 189456 119194 189512 119196
rect 189456 119142 189458 119194
rect 189458 119142 189510 119194
rect 189510 119142 189512 119194
rect 189456 119140 189512 119142
rect 189560 119194 189616 119196
rect 189560 119142 189562 119194
rect 189562 119142 189614 119194
rect 189614 119142 189616 119194
rect 189560 119140 189616 119142
rect 189664 119194 189720 119196
rect 189664 119142 189666 119194
rect 189666 119142 189718 119194
rect 189718 119142 189720 119194
rect 189664 119140 189720 119142
rect 188796 118410 188852 118412
rect 188796 118358 188798 118410
rect 188798 118358 188850 118410
rect 188850 118358 188852 118410
rect 188796 118356 188852 118358
rect 188900 118410 188956 118412
rect 188900 118358 188902 118410
rect 188902 118358 188954 118410
rect 188954 118358 188956 118410
rect 188900 118356 188956 118358
rect 189004 118410 189060 118412
rect 189004 118358 189006 118410
rect 189006 118358 189058 118410
rect 189058 118358 189060 118410
rect 189004 118356 189060 118358
rect 189456 117626 189512 117628
rect 189456 117574 189458 117626
rect 189458 117574 189510 117626
rect 189510 117574 189512 117626
rect 189456 117572 189512 117574
rect 189560 117626 189616 117628
rect 189560 117574 189562 117626
rect 189562 117574 189614 117626
rect 189614 117574 189616 117626
rect 189560 117572 189616 117574
rect 189664 117626 189720 117628
rect 189664 117574 189666 117626
rect 189666 117574 189718 117626
rect 189718 117574 189720 117626
rect 189664 117572 189720 117574
rect 188796 116842 188852 116844
rect 188796 116790 188798 116842
rect 188798 116790 188850 116842
rect 188850 116790 188852 116842
rect 188796 116788 188852 116790
rect 188900 116842 188956 116844
rect 188900 116790 188902 116842
rect 188902 116790 188954 116842
rect 188954 116790 188956 116842
rect 188900 116788 188956 116790
rect 189004 116842 189060 116844
rect 189004 116790 189006 116842
rect 189006 116790 189058 116842
rect 189058 116790 189060 116842
rect 189004 116788 189060 116790
rect 189456 116058 189512 116060
rect 189456 116006 189458 116058
rect 189458 116006 189510 116058
rect 189510 116006 189512 116058
rect 189456 116004 189512 116006
rect 189560 116058 189616 116060
rect 189560 116006 189562 116058
rect 189562 116006 189614 116058
rect 189614 116006 189616 116058
rect 189560 116004 189616 116006
rect 189664 116058 189720 116060
rect 189664 116006 189666 116058
rect 189666 116006 189718 116058
rect 189718 116006 189720 116058
rect 189664 116004 189720 116006
rect 188796 115274 188852 115276
rect 188796 115222 188798 115274
rect 188798 115222 188850 115274
rect 188850 115222 188852 115274
rect 188796 115220 188852 115222
rect 188900 115274 188956 115276
rect 188900 115222 188902 115274
rect 188902 115222 188954 115274
rect 188954 115222 188956 115274
rect 188900 115220 188956 115222
rect 189004 115274 189060 115276
rect 189004 115222 189006 115274
rect 189006 115222 189058 115274
rect 189058 115222 189060 115274
rect 189004 115220 189060 115222
rect 189456 114490 189512 114492
rect 189456 114438 189458 114490
rect 189458 114438 189510 114490
rect 189510 114438 189512 114490
rect 189456 114436 189512 114438
rect 189560 114490 189616 114492
rect 189560 114438 189562 114490
rect 189562 114438 189614 114490
rect 189614 114438 189616 114490
rect 189560 114436 189616 114438
rect 189664 114490 189720 114492
rect 189664 114438 189666 114490
rect 189666 114438 189718 114490
rect 189718 114438 189720 114490
rect 189664 114436 189720 114438
rect 188796 113706 188852 113708
rect 188796 113654 188798 113706
rect 188798 113654 188850 113706
rect 188850 113654 188852 113706
rect 188796 113652 188852 113654
rect 188900 113706 188956 113708
rect 188900 113654 188902 113706
rect 188902 113654 188954 113706
rect 188954 113654 188956 113706
rect 188900 113652 188956 113654
rect 189004 113706 189060 113708
rect 189004 113654 189006 113706
rect 189006 113654 189058 113706
rect 189058 113654 189060 113706
rect 189004 113652 189060 113654
rect 189456 112922 189512 112924
rect 189456 112870 189458 112922
rect 189458 112870 189510 112922
rect 189510 112870 189512 112922
rect 189456 112868 189512 112870
rect 189560 112922 189616 112924
rect 189560 112870 189562 112922
rect 189562 112870 189614 112922
rect 189614 112870 189616 112922
rect 189560 112868 189616 112870
rect 189664 112922 189720 112924
rect 189664 112870 189666 112922
rect 189666 112870 189718 112922
rect 189718 112870 189720 112922
rect 189664 112868 189720 112870
rect 188796 112138 188852 112140
rect 188796 112086 188798 112138
rect 188798 112086 188850 112138
rect 188850 112086 188852 112138
rect 188796 112084 188852 112086
rect 188900 112138 188956 112140
rect 188900 112086 188902 112138
rect 188902 112086 188954 112138
rect 188954 112086 188956 112138
rect 188900 112084 188956 112086
rect 189004 112138 189060 112140
rect 189004 112086 189006 112138
rect 189006 112086 189058 112138
rect 189058 112086 189060 112138
rect 189004 112084 189060 112086
rect 189456 111354 189512 111356
rect 189456 111302 189458 111354
rect 189458 111302 189510 111354
rect 189510 111302 189512 111354
rect 189456 111300 189512 111302
rect 189560 111354 189616 111356
rect 189560 111302 189562 111354
rect 189562 111302 189614 111354
rect 189614 111302 189616 111354
rect 189560 111300 189616 111302
rect 189664 111354 189720 111356
rect 189664 111302 189666 111354
rect 189666 111302 189718 111354
rect 189718 111302 189720 111354
rect 189664 111300 189720 111302
rect 188796 110570 188852 110572
rect 188796 110518 188798 110570
rect 188798 110518 188850 110570
rect 188850 110518 188852 110570
rect 188796 110516 188852 110518
rect 188900 110570 188956 110572
rect 188900 110518 188902 110570
rect 188902 110518 188954 110570
rect 188954 110518 188956 110570
rect 188900 110516 188956 110518
rect 189004 110570 189060 110572
rect 189004 110518 189006 110570
rect 189006 110518 189058 110570
rect 189058 110518 189060 110570
rect 189004 110516 189060 110518
rect 189456 109786 189512 109788
rect 189456 109734 189458 109786
rect 189458 109734 189510 109786
rect 189510 109734 189512 109786
rect 189456 109732 189512 109734
rect 189560 109786 189616 109788
rect 189560 109734 189562 109786
rect 189562 109734 189614 109786
rect 189614 109734 189616 109786
rect 189560 109732 189616 109734
rect 189664 109786 189720 109788
rect 189664 109734 189666 109786
rect 189666 109734 189718 109786
rect 189718 109734 189720 109786
rect 189664 109732 189720 109734
rect 188796 109002 188852 109004
rect 188796 108950 188798 109002
rect 188798 108950 188850 109002
rect 188850 108950 188852 109002
rect 188796 108948 188852 108950
rect 188900 109002 188956 109004
rect 188900 108950 188902 109002
rect 188902 108950 188954 109002
rect 188954 108950 188956 109002
rect 188900 108948 188956 108950
rect 189004 109002 189060 109004
rect 189004 108950 189006 109002
rect 189006 108950 189058 109002
rect 189058 108950 189060 109002
rect 189004 108948 189060 108950
rect 189456 108218 189512 108220
rect 189456 108166 189458 108218
rect 189458 108166 189510 108218
rect 189510 108166 189512 108218
rect 189456 108164 189512 108166
rect 189560 108218 189616 108220
rect 189560 108166 189562 108218
rect 189562 108166 189614 108218
rect 189614 108166 189616 108218
rect 189560 108164 189616 108166
rect 189664 108218 189720 108220
rect 189664 108166 189666 108218
rect 189666 108166 189718 108218
rect 189718 108166 189720 108218
rect 189664 108164 189720 108166
rect 188796 107434 188852 107436
rect 188796 107382 188798 107434
rect 188798 107382 188850 107434
rect 188850 107382 188852 107434
rect 188796 107380 188852 107382
rect 188900 107434 188956 107436
rect 188900 107382 188902 107434
rect 188902 107382 188954 107434
rect 188954 107382 188956 107434
rect 188900 107380 188956 107382
rect 189004 107434 189060 107436
rect 189004 107382 189006 107434
rect 189006 107382 189058 107434
rect 189058 107382 189060 107434
rect 189004 107380 189060 107382
rect 189456 106650 189512 106652
rect 189456 106598 189458 106650
rect 189458 106598 189510 106650
rect 189510 106598 189512 106650
rect 189456 106596 189512 106598
rect 189560 106650 189616 106652
rect 189560 106598 189562 106650
rect 189562 106598 189614 106650
rect 189614 106598 189616 106650
rect 189560 106596 189616 106598
rect 189664 106650 189720 106652
rect 189664 106598 189666 106650
rect 189666 106598 189718 106650
rect 189718 106598 189720 106650
rect 189664 106596 189720 106598
rect 188796 105866 188852 105868
rect 188796 105814 188798 105866
rect 188798 105814 188850 105866
rect 188850 105814 188852 105866
rect 188796 105812 188852 105814
rect 188900 105866 188956 105868
rect 188900 105814 188902 105866
rect 188902 105814 188954 105866
rect 188954 105814 188956 105866
rect 188900 105812 188956 105814
rect 189004 105866 189060 105868
rect 189004 105814 189006 105866
rect 189006 105814 189058 105866
rect 189058 105814 189060 105866
rect 189004 105812 189060 105814
rect 189456 105082 189512 105084
rect 189456 105030 189458 105082
rect 189458 105030 189510 105082
rect 189510 105030 189512 105082
rect 189456 105028 189512 105030
rect 189560 105082 189616 105084
rect 189560 105030 189562 105082
rect 189562 105030 189614 105082
rect 189614 105030 189616 105082
rect 189560 105028 189616 105030
rect 189664 105082 189720 105084
rect 189664 105030 189666 105082
rect 189666 105030 189718 105082
rect 189718 105030 189720 105082
rect 189664 105028 189720 105030
rect 188796 104298 188852 104300
rect 188796 104246 188798 104298
rect 188798 104246 188850 104298
rect 188850 104246 188852 104298
rect 188796 104244 188852 104246
rect 188900 104298 188956 104300
rect 188900 104246 188902 104298
rect 188902 104246 188954 104298
rect 188954 104246 188956 104298
rect 188900 104244 188956 104246
rect 189004 104298 189060 104300
rect 189004 104246 189006 104298
rect 189006 104246 189058 104298
rect 189058 104246 189060 104298
rect 189004 104244 189060 104246
rect 189456 103514 189512 103516
rect 189456 103462 189458 103514
rect 189458 103462 189510 103514
rect 189510 103462 189512 103514
rect 189456 103460 189512 103462
rect 189560 103514 189616 103516
rect 189560 103462 189562 103514
rect 189562 103462 189614 103514
rect 189614 103462 189616 103514
rect 189560 103460 189616 103462
rect 189664 103514 189720 103516
rect 189664 103462 189666 103514
rect 189666 103462 189718 103514
rect 189718 103462 189720 103514
rect 189664 103460 189720 103462
rect 188796 102730 188852 102732
rect 188796 102678 188798 102730
rect 188798 102678 188850 102730
rect 188850 102678 188852 102730
rect 188796 102676 188852 102678
rect 188900 102730 188956 102732
rect 188900 102678 188902 102730
rect 188902 102678 188954 102730
rect 188954 102678 188956 102730
rect 188900 102676 188956 102678
rect 189004 102730 189060 102732
rect 189004 102678 189006 102730
rect 189006 102678 189058 102730
rect 189058 102678 189060 102730
rect 189004 102676 189060 102678
rect 189456 101946 189512 101948
rect 189456 101894 189458 101946
rect 189458 101894 189510 101946
rect 189510 101894 189512 101946
rect 189456 101892 189512 101894
rect 189560 101946 189616 101948
rect 189560 101894 189562 101946
rect 189562 101894 189614 101946
rect 189614 101894 189616 101946
rect 189560 101892 189616 101894
rect 189664 101946 189720 101948
rect 189664 101894 189666 101946
rect 189666 101894 189718 101946
rect 189718 101894 189720 101946
rect 189664 101892 189720 101894
rect 188796 101162 188852 101164
rect 188796 101110 188798 101162
rect 188798 101110 188850 101162
rect 188850 101110 188852 101162
rect 188796 101108 188852 101110
rect 188900 101162 188956 101164
rect 188900 101110 188902 101162
rect 188902 101110 188954 101162
rect 188954 101110 188956 101162
rect 188900 101108 188956 101110
rect 189004 101162 189060 101164
rect 189004 101110 189006 101162
rect 189006 101110 189058 101162
rect 189058 101110 189060 101162
rect 189004 101108 189060 101110
rect 189456 100378 189512 100380
rect 189456 100326 189458 100378
rect 189458 100326 189510 100378
rect 189510 100326 189512 100378
rect 189456 100324 189512 100326
rect 189560 100378 189616 100380
rect 189560 100326 189562 100378
rect 189562 100326 189614 100378
rect 189614 100326 189616 100378
rect 189560 100324 189616 100326
rect 189664 100378 189720 100380
rect 189664 100326 189666 100378
rect 189666 100326 189718 100378
rect 189718 100326 189720 100378
rect 189664 100324 189720 100326
rect 188796 99594 188852 99596
rect 188796 99542 188798 99594
rect 188798 99542 188850 99594
rect 188850 99542 188852 99594
rect 188796 99540 188852 99542
rect 188900 99594 188956 99596
rect 188900 99542 188902 99594
rect 188902 99542 188954 99594
rect 188954 99542 188956 99594
rect 188900 99540 188956 99542
rect 189004 99594 189060 99596
rect 189004 99542 189006 99594
rect 189006 99542 189058 99594
rect 189058 99542 189060 99594
rect 189004 99540 189060 99542
rect 189456 98810 189512 98812
rect 189456 98758 189458 98810
rect 189458 98758 189510 98810
rect 189510 98758 189512 98810
rect 189456 98756 189512 98758
rect 189560 98810 189616 98812
rect 189560 98758 189562 98810
rect 189562 98758 189614 98810
rect 189614 98758 189616 98810
rect 189560 98756 189616 98758
rect 189664 98810 189720 98812
rect 189664 98758 189666 98810
rect 189666 98758 189718 98810
rect 189718 98758 189720 98810
rect 189664 98756 189720 98758
rect 188796 98026 188852 98028
rect 188796 97974 188798 98026
rect 188798 97974 188850 98026
rect 188850 97974 188852 98026
rect 188796 97972 188852 97974
rect 188900 98026 188956 98028
rect 188900 97974 188902 98026
rect 188902 97974 188954 98026
rect 188954 97974 188956 98026
rect 188900 97972 188956 97974
rect 189004 98026 189060 98028
rect 189004 97974 189006 98026
rect 189006 97974 189058 98026
rect 189058 97974 189060 98026
rect 189004 97972 189060 97974
rect 189456 97242 189512 97244
rect 189456 97190 189458 97242
rect 189458 97190 189510 97242
rect 189510 97190 189512 97242
rect 189456 97188 189512 97190
rect 189560 97242 189616 97244
rect 189560 97190 189562 97242
rect 189562 97190 189614 97242
rect 189614 97190 189616 97242
rect 189560 97188 189616 97190
rect 189664 97242 189720 97244
rect 189664 97190 189666 97242
rect 189666 97190 189718 97242
rect 189718 97190 189720 97242
rect 189664 97188 189720 97190
rect 188796 96458 188852 96460
rect 188796 96406 188798 96458
rect 188798 96406 188850 96458
rect 188850 96406 188852 96458
rect 188796 96404 188852 96406
rect 188900 96458 188956 96460
rect 188900 96406 188902 96458
rect 188902 96406 188954 96458
rect 188954 96406 188956 96458
rect 188900 96404 188956 96406
rect 189004 96458 189060 96460
rect 189004 96406 189006 96458
rect 189006 96406 189058 96458
rect 189058 96406 189060 96458
rect 189004 96404 189060 96406
rect 189456 95674 189512 95676
rect 189456 95622 189458 95674
rect 189458 95622 189510 95674
rect 189510 95622 189512 95674
rect 189456 95620 189512 95622
rect 189560 95674 189616 95676
rect 189560 95622 189562 95674
rect 189562 95622 189614 95674
rect 189614 95622 189616 95674
rect 189560 95620 189616 95622
rect 189664 95674 189720 95676
rect 189664 95622 189666 95674
rect 189666 95622 189718 95674
rect 189718 95622 189720 95674
rect 189664 95620 189720 95622
rect 188796 94890 188852 94892
rect 188796 94838 188798 94890
rect 188798 94838 188850 94890
rect 188850 94838 188852 94890
rect 188796 94836 188852 94838
rect 188900 94890 188956 94892
rect 188900 94838 188902 94890
rect 188902 94838 188954 94890
rect 188954 94838 188956 94890
rect 188900 94836 188956 94838
rect 189004 94890 189060 94892
rect 189004 94838 189006 94890
rect 189006 94838 189058 94890
rect 189058 94838 189060 94890
rect 189004 94836 189060 94838
rect 189456 94106 189512 94108
rect 189456 94054 189458 94106
rect 189458 94054 189510 94106
rect 189510 94054 189512 94106
rect 189456 94052 189512 94054
rect 189560 94106 189616 94108
rect 189560 94054 189562 94106
rect 189562 94054 189614 94106
rect 189614 94054 189616 94106
rect 189560 94052 189616 94054
rect 189664 94106 189720 94108
rect 189664 94054 189666 94106
rect 189666 94054 189718 94106
rect 189718 94054 189720 94106
rect 189664 94052 189720 94054
rect 190652 93660 190708 93716
rect 188796 93322 188852 93324
rect 188796 93270 188798 93322
rect 188798 93270 188850 93322
rect 188850 93270 188852 93322
rect 188796 93268 188852 93270
rect 188900 93322 188956 93324
rect 188900 93270 188902 93322
rect 188902 93270 188954 93322
rect 188954 93270 188956 93322
rect 188900 93268 188956 93270
rect 189004 93322 189060 93324
rect 189004 93270 189006 93322
rect 189006 93270 189058 93322
rect 189058 93270 189060 93322
rect 189004 93268 189060 93270
rect 189456 92538 189512 92540
rect 189456 92486 189458 92538
rect 189458 92486 189510 92538
rect 189510 92486 189512 92538
rect 189456 92484 189512 92486
rect 189560 92538 189616 92540
rect 189560 92486 189562 92538
rect 189562 92486 189614 92538
rect 189614 92486 189616 92538
rect 189560 92484 189616 92486
rect 189664 92538 189720 92540
rect 189664 92486 189666 92538
rect 189666 92486 189718 92538
rect 189718 92486 189720 92538
rect 189664 92484 189720 92486
rect 188796 91754 188852 91756
rect 188796 91702 188798 91754
rect 188798 91702 188850 91754
rect 188850 91702 188852 91754
rect 188796 91700 188852 91702
rect 188900 91754 188956 91756
rect 188900 91702 188902 91754
rect 188902 91702 188954 91754
rect 188954 91702 188956 91754
rect 188900 91700 188956 91702
rect 189004 91754 189060 91756
rect 189004 91702 189006 91754
rect 189006 91702 189058 91754
rect 189058 91702 189060 91754
rect 189004 91700 189060 91702
rect 189456 90970 189512 90972
rect 189456 90918 189458 90970
rect 189458 90918 189510 90970
rect 189510 90918 189512 90970
rect 189456 90916 189512 90918
rect 189560 90970 189616 90972
rect 189560 90918 189562 90970
rect 189562 90918 189614 90970
rect 189614 90918 189616 90970
rect 189560 90916 189616 90918
rect 189664 90970 189720 90972
rect 189664 90918 189666 90970
rect 189666 90918 189718 90970
rect 189718 90918 189720 90970
rect 189664 90916 189720 90918
rect 188796 90186 188852 90188
rect 188796 90134 188798 90186
rect 188798 90134 188850 90186
rect 188850 90134 188852 90186
rect 188796 90132 188852 90134
rect 188900 90186 188956 90188
rect 188900 90134 188902 90186
rect 188902 90134 188954 90186
rect 188954 90134 188956 90186
rect 188900 90132 188956 90134
rect 189004 90186 189060 90188
rect 189004 90134 189006 90186
rect 189006 90134 189058 90186
rect 189058 90134 189060 90186
rect 189004 90132 189060 90134
rect 189456 89402 189512 89404
rect 189456 89350 189458 89402
rect 189458 89350 189510 89402
rect 189510 89350 189512 89402
rect 189456 89348 189512 89350
rect 189560 89402 189616 89404
rect 189560 89350 189562 89402
rect 189562 89350 189614 89402
rect 189614 89350 189616 89402
rect 189560 89348 189616 89350
rect 189664 89402 189720 89404
rect 189664 89350 189666 89402
rect 189666 89350 189718 89402
rect 189718 89350 189720 89402
rect 189664 89348 189720 89350
rect 188796 88618 188852 88620
rect 188796 88566 188798 88618
rect 188798 88566 188850 88618
rect 188850 88566 188852 88618
rect 188796 88564 188852 88566
rect 188900 88618 188956 88620
rect 188900 88566 188902 88618
rect 188902 88566 188954 88618
rect 188954 88566 188956 88618
rect 188900 88564 188956 88566
rect 189004 88618 189060 88620
rect 189004 88566 189006 88618
rect 189006 88566 189058 88618
rect 189058 88566 189060 88618
rect 189004 88564 189060 88566
rect 189456 87834 189512 87836
rect 189456 87782 189458 87834
rect 189458 87782 189510 87834
rect 189510 87782 189512 87834
rect 189456 87780 189512 87782
rect 189560 87834 189616 87836
rect 189560 87782 189562 87834
rect 189562 87782 189614 87834
rect 189614 87782 189616 87834
rect 189560 87780 189616 87782
rect 189664 87834 189720 87836
rect 189664 87782 189666 87834
rect 189666 87782 189718 87834
rect 189718 87782 189720 87834
rect 189664 87780 189720 87782
rect 188796 87050 188852 87052
rect 188796 86998 188798 87050
rect 188798 86998 188850 87050
rect 188850 86998 188852 87050
rect 188796 86996 188852 86998
rect 188900 87050 188956 87052
rect 188900 86998 188902 87050
rect 188902 86998 188954 87050
rect 188954 86998 188956 87050
rect 188900 86996 188956 86998
rect 189004 87050 189060 87052
rect 189004 86998 189006 87050
rect 189006 86998 189058 87050
rect 189058 86998 189060 87050
rect 189004 86996 189060 86998
rect 189456 86266 189512 86268
rect 189456 86214 189458 86266
rect 189458 86214 189510 86266
rect 189510 86214 189512 86266
rect 189456 86212 189512 86214
rect 189560 86266 189616 86268
rect 189560 86214 189562 86266
rect 189562 86214 189614 86266
rect 189614 86214 189616 86266
rect 189560 86212 189616 86214
rect 189664 86266 189720 86268
rect 189664 86214 189666 86266
rect 189666 86214 189718 86266
rect 189718 86214 189720 86266
rect 189664 86212 189720 86214
rect 188796 85482 188852 85484
rect 188796 85430 188798 85482
rect 188798 85430 188850 85482
rect 188850 85430 188852 85482
rect 188796 85428 188852 85430
rect 188900 85482 188956 85484
rect 188900 85430 188902 85482
rect 188902 85430 188954 85482
rect 188954 85430 188956 85482
rect 188900 85428 188956 85430
rect 189004 85482 189060 85484
rect 189004 85430 189006 85482
rect 189006 85430 189058 85482
rect 189058 85430 189060 85482
rect 189004 85428 189060 85430
rect 189456 84698 189512 84700
rect 189456 84646 189458 84698
rect 189458 84646 189510 84698
rect 189510 84646 189512 84698
rect 189456 84644 189512 84646
rect 189560 84698 189616 84700
rect 189560 84646 189562 84698
rect 189562 84646 189614 84698
rect 189614 84646 189616 84698
rect 189560 84644 189616 84646
rect 189664 84698 189720 84700
rect 189664 84646 189666 84698
rect 189666 84646 189718 84698
rect 189718 84646 189720 84698
rect 189664 84644 189720 84646
rect 188796 83914 188852 83916
rect 188796 83862 188798 83914
rect 188798 83862 188850 83914
rect 188850 83862 188852 83914
rect 188796 83860 188852 83862
rect 188900 83914 188956 83916
rect 188900 83862 188902 83914
rect 188902 83862 188954 83914
rect 188954 83862 188956 83914
rect 188900 83860 188956 83862
rect 189004 83914 189060 83916
rect 189004 83862 189006 83914
rect 189006 83862 189058 83914
rect 189058 83862 189060 83914
rect 189004 83860 189060 83862
rect 189456 83130 189512 83132
rect 189456 83078 189458 83130
rect 189458 83078 189510 83130
rect 189510 83078 189512 83130
rect 189456 83076 189512 83078
rect 189560 83130 189616 83132
rect 189560 83078 189562 83130
rect 189562 83078 189614 83130
rect 189614 83078 189616 83130
rect 189560 83076 189616 83078
rect 189664 83130 189720 83132
rect 189664 83078 189666 83130
rect 189666 83078 189718 83130
rect 189718 83078 189720 83130
rect 189664 83076 189720 83078
rect 188796 82346 188852 82348
rect 188796 82294 188798 82346
rect 188798 82294 188850 82346
rect 188850 82294 188852 82346
rect 188796 82292 188852 82294
rect 188900 82346 188956 82348
rect 188900 82294 188902 82346
rect 188902 82294 188954 82346
rect 188954 82294 188956 82346
rect 188900 82292 188956 82294
rect 189004 82346 189060 82348
rect 189004 82294 189006 82346
rect 189006 82294 189058 82346
rect 189058 82294 189060 82346
rect 189004 82292 189060 82294
rect 189456 81562 189512 81564
rect 189456 81510 189458 81562
rect 189458 81510 189510 81562
rect 189510 81510 189512 81562
rect 189456 81508 189512 81510
rect 189560 81562 189616 81564
rect 189560 81510 189562 81562
rect 189562 81510 189614 81562
rect 189614 81510 189616 81562
rect 189560 81508 189616 81510
rect 189664 81562 189720 81564
rect 189664 81510 189666 81562
rect 189666 81510 189718 81562
rect 189718 81510 189720 81562
rect 189664 81508 189720 81510
rect 188796 80778 188852 80780
rect 188796 80726 188798 80778
rect 188798 80726 188850 80778
rect 188850 80726 188852 80778
rect 188796 80724 188852 80726
rect 188900 80778 188956 80780
rect 188900 80726 188902 80778
rect 188902 80726 188954 80778
rect 188954 80726 188956 80778
rect 188900 80724 188956 80726
rect 189004 80778 189060 80780
rect 189004 80726 189006 80778
rect 189006 80726 189058 80778
rect 189058 80726 189060 80778
rect 189004 80724 189060 80726
rect 189456 79994 189512 79996
rect 189456 79942 189458 79994
rect 189458 79942 189510 79994
rect 189510 79942 189512 79994
rect 189456 79940 189512 79942
rect 189560 79994 189616 79996
rect 189560 79942 189562 79994
rect 189562 79942 189614 79994
rect 189614 79942 189616 79994
rect 189560 79940 189616 79942
rect 189664 79994 189720 79996
rect 189664 79942 189666 79994
rect 189666 79942 189718 79994
rect 189718 79942 189720 79994
rect 189664 79940 189720 79942
rect 188796 79210 188852 79212
rect 188796 79158 188798 79210
rect 188798 79158 188850 79210
rect 188850 79158 188852 79210
rect 188796 79156 188852 79158
rect 188900 79210 188956 79212
rect 188900 79158 188902 79210
rect 188902 79158 188954 79210
rect 188954 79158 188956 79210
rect 188900 79156 188956 79158
rect 189004 79210 189060 79212
rect 189004 79158 189006 79210
rect 189006 79158 189058 79210
rect 189058 79158 189060 79210
rect 189004 79156 189060 79158
rect 189456 78426 189512 78428
rect 189456 78374 189458 78426
rect 189458 78374 189510 78426
rect 189510 78374 189512 78426
rect 189456 78372 189512 78374
rect 189560 78426 189616 78428
rect 189560 78374 189562 78426
rect 189562 78374 189614 78426
rect 189614 78374 189616 78426
rect 189560 78372 189616 78374
rect 189664 78426 189720 78428
rect 189664 78374 189666 78426
rect 189666 78374 189718 78426
rect 189718 78374 189720 78426
rect 189664 78372 189720 78374
rect 188796 77642 188852 77644
rect 188796 77590 188798 77642
rect 188798 77590 188850 77642
rect 188850 77590 188852 77642
rect 188796 77588 188852 77590
rect 188900 77642 188956 77644
rect 188900 77590 188902 77642
rect 188902 77590 188954 77642
rect 188954 77590 188956 77642
rect 188900 77588 188956 77590
rect 189004 77642 189060 77644
rect 189004 77590 189006 77642
rect 189006 77590 189058 77642
rect 189058 77590 189060 77642
rect 189004 77588 189060 77590
rect 189456 76858 189512 76860
rect 189456 76806 189458 76858
rect 189458 76806 189510 76858
rect 189510 76806 189512 76858
rect 189456 76804 189512 76806
rect 189560 76858 189616 76860
rect 189560 76806 189562 76858
rect 189562 76806 189614 76858
rect 189614 76806 189616 76858
rect 189560 76804 189616 76806
rect 189664 76858 189720 76860
rect 189664 76806 189666 76858
rect 189666 76806 189718 76858
rect 189718 76806 189720 76858
rect 189664 76804 189720 76806
rect 188796 76074 188852 76076
rect 188796 76022 188798 76074
rect 188798 76022 188850 76074
rect 188850 76022 188852 76074
rect 188796 76020 188852 76022
rect 188900 76074 188956 76076
rect 188900 76022 188902 76074
rect 188902 76022 188954 76074
rect 188954 76022 188956 76074
rect 188900 76020 188956 76022
rect 189004 76074 189060 76076
rect 189004 76022 189006 76074
rect 189006 76022 189058 76074
rect 189058 76022 189060 76074
rect 189004 76020 189060 76022
rect 189456 75290 189512 75292
rect 189456 75238 189458 75290
rect 189458 75238 189510 75290
rect 189510 75238 189512 75290
rect 189456 75236 189512 75238
rect 189560 75290 189616 75292
rect 189560 75238 189562 75290
rect 189562 75238 189614 75290
rect 189614 75238 189616 75290
rect 189560 75236 189616 75238
rect 189664 75290 189720 75292
rect 189664 75238 189666 75290
rect 189666 75238 189718 75290
rect 189718 75238 189720 75290
rect 189664 75236 189720 75238
rect 188796 74506 188852 74508
rect 188796 74454 188798 74506
rect 188798 74454 188850 74506
rect 188850 74454 188852 74506
rect 188796 74452 188852 74454
rect 188900 74506 188956 74508
rect 188900 74454 188902 74506
rect 188902 74454 188954 74506
rect 188954 74454 188956 74506
rect 188900 74452 188956 74454
rect 189004 74506 189060 74508
rect 189004 74454 189006 74506
rect 189006 74454 189058 74506
rect 189058 74454 189060 74506
rect 189004 74452 189060 74454
rect 189456 73722 189512 73724
rect 189456 73670 189458 73722
rect 189458 73670 189510 73722
rect 189510 73670 189512 73722
rect 189456 73668 189512 73670
rect 189560 73722 189616 73724
rect 189560 73670 189562 73722
rect 189562 73670 189614 73722
rect 189614 73670 189616 73722
rect 189560 73668 189616 73670
rect 189664 73722 189720 73724
rect 189664 73670 189666 73722
rect 189666 73670 189718 73722
rect 189718 73670 189720 73722
rect 189664 73668 189720 73670
rect 188796 72938 188852 72940
rect 188796 72886 188798 72938
rect 188798 72886 188850 72938
rect 188850 72886 188852 72938
rect 188796 72884 188852 72886
rect 188900 72938 188956 72940
rect 188900 72886 188902 72938
rect 188902 72886 188954 72938
rect 188954 72886 188956 72938
rect 188900 72884 188956 72886
rect 189004 72938 189060 72940
rect 189004 72886 189006 72938
rect 189006 72886 189058 72938
rect 189058 72886 189060 72938
rect 189004 72884 189060 72886
rect 189456 72154 189512 72156
rect 189456 72102 189458 72154
rect 189458 72102 189510 72154
rect 189510 72102 189512 72154
rect 189456 72100 189512 72102
rect 189560 72154 189616 72156
rect 189560 72102 189562 72154
rect 189562 72102 189614 72154
rect 189614 72102 189616 72154
rect 189560 72100 189616 72102
rect 189664 72154 189720 72156
rect 189664 72102 189666 72154
rect 189666 72102 189718 72154
rect 189718 72102 189720 72154
rect 189664 72100 189720 72102
rect 188796 71370 188852 71372
rect 188796 71318 188798 71370
rect 188798 71318 188850 71370
rect 188850 71318 188852 71370
rect 188796 71316 188852 71318
rect 188900 71370 188956 71372
rect 188900 71318 188902 71370
rect 188902 71318 188954 71370
rect 188954 71318 188956 71370
rect 188900 71316 188956 71318
rect 189004 71370 189060 71372
rect 189004 71318 189006 71370
rect 189006 71318 189058 71370
rect 189058 71318 189060 71370
rect 189004 71316 189060 71318
rect 189456 70586 189512 70588
rect 189456 70534 189458 70586
rect 189458 70534 189510 70586
rect 189510 70534 189512 70586
rect 189456 70532 189512 70534
rect 189560 70586 189616 70588
rect 189560 70534 189562 70586
rect 189562 70534 189614 70586
rect 189614 70534 189616 70586
rect 189560 70532 189616 70534
rect 189664 70586 189720 70588
rect 189664 70534 189666 70586
rect 189666 70534 189718 70586
rect 189718 70534 189720 70586
rect 189664 70532 189720 70534
rect 188796 69802 188852 69804
rect 188796 69750 188798 69802
rect 188798 69750 188850 69802
rect 188850 69750 188852 69802
rect 188796 69748 188852 69750
rect 188900 69802 188956 69804
rect 188900 69750 188902 69802
rect 188902 69750 188954 69802
rect 188954 69750 188956 69802
rect 188900 69748 188956 69750
rect 189004 69802 189060 69804
rect 189004 69750 189006 69802
rect 189006 69750 189058 69802
rect 189058 69750 189060 69802
rect 189004 69748 189060 69750
rect 189456 69018 189512 69020
rect 189456 68966 189458 69018
rect 189458 68966 189510 69018
rect 189510 68966 189512 69018
rect 189456 68964 189512 68966
rect 189560 69018 189616 69020
rect 189560 68966 189562 69018
rect 189562 68966 189614 69018
rect 189614 68966 189616 69018
rect 189560 68964 189616 68966
rect 189664 69018 189720 69020
rect 189664 68966 189666 69018
rect 189666 68966 189718 69018
rect 189718 68966 189720 69018
rect 189664 68964 189720 68966
rect 188796 68234 188852 68236
rect 188796 68182 188798 68234
rect 188798 68182 188850 68234
rect 188850 68182 188852 68234
rect 188796 68180 188852 68182
rect 188900 68234 188956 68236
rect 188900 68182 188902 68234
rect 188902 68182 188954 68234
rect 188954 68182 188956 68234
rect 188900 68180 188956 68182
rect 189004 68234 189060 68236
rect 189004 68182 189006 68234
rect 189006 68182 189058 68234
rect 189058 68182 189060 68234
rect 189004 68180 189060 68182
rect 189456 67450 189512 67452
rect 189456 67398 189458 67450
rect 189458 67398 189510 67450
rect 189510 67398 189512 67450
rect 189456 67396 189512 67398
rect 189560 67450 189616 67452
rect 189560 67398 189562 67450
rect 189562 67398 189614 67450
rect 189614 67398 189616 67450
rect 189560 67396 189616 67398
rect 189664 67450 189720 67452
rect 189664 67398 189666 67450
rect 189666 67398 189718 67450
rect 189718 67398 189720 67450
rect 189664 67396 189720 67398
rect 187292 67004 187348 67060
rect 173964 38668 174020 38724
rect 156380 37996 156436 38052
rect 85148 31836 85204 31892
rect 75516 21756 75572 21812
rect 75628 29372 75684 29428
rect 154588 29372 154644 29428
rect 149548 26124 149604 26180
rect 78876 25452 78932 25508
rect 149548 22876 149604 22932
rect 78876 22652 78932 22708
rect 97132 22652 97188 22708
rect 82908 21196 82964 21252
rect 75628 20412 75684 20468
rect 82460 20412 82516 20468
rect 78988 17106 79044 17108
rect 78988 17054 78990 17106
rect 78990 17054 79042 17106
rect 79042 17054 79044 17106
rect 78988 17052 79044 17054
rect 140028 22652 140084 22708
rect 111244 21084 111300 21140
rect 97296 17274 97352 17276
rect 97296 17222 97298 17274
rect 97298 17222 97350 17274
rect 97350 17222 97352 17274
rect 97296 17220 97352 17222
rect 97400 17274 97456 17276
rect 97400 17222 97402 17274
rect 97402 17222 97454 17274
rect 97454 17222 97456 17274
rect 97400 17220 97456 17222
rect 97504 17274 97560 17276
rect 97504 17222 97506 17274
rect 97506 17222 97558 17274
rect 97558 17222 97560 17274
rect 97504 17220 97560 17222
rect 128016 17274 128072 17276
rect 128016 17222 128018 17274
rect 128018 17222 128070 17274
rect 128070 17222 128072 17274
rect 128016 17220 128072 17222
rect 128120 17274 128176 17276
rect 128120 17222 128122 17274
rect 128122 17222 128174 17274
rect 128174 17222 128176 17274
rect 128120 17220 128176 17222
rect 128224 17274 128280 17276
rect 128224 17222 128226 17274
rect 128226 17222 128278 17274
rect 128278 17222 128280 17274
rect 128224 17220 128280 17222
rect 188796 66666 188852 66668
rect 188796 66614 188798 66666
rect 188798 66614 188850 66666
rect 188850 66614 188852 66666
rect 188796 66612 188852 66614
rect 188900 66666 188956 66668
rect 188900 66614 188902 66666
rect 188902 66614 188954 66666
rect 188954 66614 188956 66666
rect 188900 66612 188956 66614
rect 189004 66666 189060 66668
rect 189004 66614 189006 66666
rect 189006 66614 189058 66666
rect 189058 66614 189060 66666
rect 189004 66612 189060 66614
rect 189456 65882 189512 65884
rect 189456 65830 189458 65882
rect 189458 65830 189510 65882
rect 189510 65830 189512 65882
rect 189456 65828 189512 65830
rect 189560 65882 189616 65884
rect 189560 65830 189562 65882
rect 189562 65830 189614 65882
rect 189614 65830 189616 65882
rect 189560 65828 189616 65830
rect 189664 65882 189720 65884
rect 189664 65830 189666 65882
rect 189666 65830 189718 65882
rect 189718 65830 189720 65882
rect 189664 65828 189720 65830
rect 188796 65098 188852 65100
rect 188796 65046 188798 65098
rect 188798 65046 188850 65098
rect 188850 65046 188852 65098
rect 188796 65044 188852 65046
rect 188900 65098 188956 65100
rect 188900 65046 188902 65098
rect 188902 65046 188954 65098
rect 188954 65046 188956 65098
rect 188900 65044 188956 65046
rect 189004 65098 189060 65100
rect 189004 65046 189006 65098
rect 189006 65046 189058 65098
rect 189058 65046 189060 65098
rect 189004 65044 189060 65046
rect 189456 64314 189512 64316
rect 189456 64262 189458 64314
rect 189458 64262 189510 64314
rect 189510 64262 189512 64314
rect 189456 64260 189512 64262
rect 189560 64314 189616 64316
rect 189560 64262 189562 64314
rect 189562 64262 189614 64314
rect 189614 64262 189616 64314
rect 189560 64260 189616 64262
rect 189664 64314 189720 64316
rect 189664 64262 189666 64314
rect 189666 64262 189718 64314
rect 189718 64262 189720 64314
rect 189664 64260 189720 64262
rect 188796 63530 188852 63532
rect 188796 63478 188798 63530
rect 188798 63478 188850 63530
rect 188850 63478 188852 63530
rect 188796 63476 188852 63478
rect 188900 63530 188956 63532
rect 188900 63478 188902 63530
rect 188902 63478 188954 63530
rect 188954 63478 188956 63530
rect 188900 63476 188956 63478
rect 189004 63530 189060 63532
rect 189004 63478 189006 63530
rect 189006 63478 189058 63530
rect 189058 63478 189060 63530
rect 189004 63476 189060 63478
rect 189456 62746 189512 62748
rect 189456 62694 189458 62746
rect 189458 62694 189510 62746
rect 189510 62694 189512 62746
rect 189456 62692 189512 62694
rect 189560 62746 189616 62748
rect 189560 62694 189562 62746
rect 189562 62694 189614 62746
rect 189614 62694 189616 62746
rect 189560 62692 189616 62694
rect 189664 62746 189720 62748
rect 189664 62694 189666 62746
rect 189666 62694 189718 62746
rect 189718 62694 189720 62746
rect 189664 62692 189720 62694
rect 188796 61962 188852 61964
rect 188796 61910 188798 61962
rect 188798 61910 188850 61962
rect 188850 61910 188852 61962
rect 188796 61908 188852 61910
rect 188900 61962 188956 61964
rect 188900 61910 188902 61962
rect 188902 61910 188954 61962
rect 188954 61910 188956 61962
rect 188900 61908 188956 61910
rect 189004 61962 189060 61964
rect 189004 61910 189006 61962
rect 189006 61910 189058 61962
rect 189058 61910 189060 61962
rect 189004 61908 189060 61910
rect 189456 61178 189512 61180
rect 189456 61126 189458 61178
rect 189458 61126 189510 61178
rect 189510 61126 189512 61178
rect 189456 61124 189512 61126
rect 189560 61178 189616 61180
rect 189560 61126 189562 61178
rect 189562 61126 189614 61178
rect 189614 61126 189616 61178
rect 189560 61124 189616 61126
rect 189664 61178 189720 61180
rect 189664 61126 189666 61178
rect 189666 61126 189718 61178
rect 189718 61126 189720 61178
rect 189664 61124 189720 61126
rect 188796 60394 188852 60396
rect 188796 60342 188798 60394
rect 188798 60342 188850 60394
rect 188850 60342 188852 60394
rect 188796 60340 188852 60342
rect 188900 60394 188956 60396
rect 188900 60342 188902 60394
rect 188902 60342 188954 60394
rect 188954 60342 188956 60394
rect 188900 60340 188956 60342
rect 189004 60394 189060 60396
rect 189004 60342 189006 60394
rect 189006 60342 189058 60394
rect 189058 60342 189060 60394
rect 189004 60340 189060 60342
rect 189456 59610 189512 59612
rect 189456 59558 189458 59610
rect 189458 59558 189510 59610
rect 189510 59558 189512 59610
rect 189456 59556 189512 59558
rect 189560 59610 189616 59612
rect 189560 59558 189562 59610
rect 189562 59558 189614 59610
rect 189614 59558 189616 59610
rect 189560 59556 189616 59558
rect 189664 59610 189720 59612
rect 189664 59558 189666 59610
rect 189666 59558 189718 59610
rect 189718 59558 189720 59610
rect 189664 59556 189720 59558
rect 188796 58826 188852 58828
rect 188796 58774 188798 58826
rect 188798 58774 188850 58826
rect 188850 58774 188852 58826
rect 188796 58772 188852 58774
rect 188900 58826 188956 58828
rect 188900 58774 188902 58826
rect 188902 58774 188954 58826
rect 188954 58774 188956 58826
rect 188900 58772 188956 58774
rect 189004 58826 189060 58828
rect 189004 58774 189006 58826
rect 189006 58774 189058 58826
rect 189058 58774 189060 58826
rect 189004 58772 189060 58774
rect 189456 58042 189512 58044
rect 189456 57990 189458 58042
rect 189458 57990 189510 58042
rect 189510 57990 189512 58042
rect 189456 57988 189512 57990
rect 189560 58042 189616 58044
rect 189560 57990 189562 58042
rect 189562 57990 189614 58042
rect 189614 57990 189616 58042
rect 189560 57988 189616 57990
rect 189664 58042 189720 58044
rect 189664 57990 189666 58042
rect 189666 57990 189718 58042
rect 189718 57990 189720 58042
rect 189664 57988 189720 57990
rect 188796 57258 188852 57260
rect 188796 57206 188798 57258
rect 188798 57206 188850 57258
rect 188850 57206 188852 57258
rect 188796 57204 188852 57206
rect 188900 57258 188956 57260
rect 188900 57206 188902 57258
rect 188902 57206 188954 57258
rect 188954 57206 188956 57258
rect 188900 57204 188956 57206
rect 189004 57258 189060 57260
rect 189004 57206 189006 57258
rect 189006 57206 189058 57258
rect 189058 57206 189060 57258
rect 189004 57204 189060 57206
rect 189456 56474 189512 56476
rect 189456 56422 189458 56474
rect 189458 56422 189510 56474
rect 189510 56422 189512 56474
rect 189456 56420 189512 56422
rect 189560 56474 189616 56476
rect 189560 56422 189562 56474
rect 189562 56422 189614 56474
rect 189614 56422 189616 56474
rect 189560 56420 189616 56422
rect 189664 56474 189720 56476
rect 189664 56422 189666 56474
rect 189666 56422 189718 56474
rect 189718 56422 189720 56474
rect 189664 56420 189720 56422
rect 188796 55690 188852 55692
rect 188796 55638 188798 55690
rect 188798 55638 188850 55690
rect 188850 55638 188852 55690
rect 188796 55636 188852 55638
rect 188900 55690 188956 55692
rect 188900 55638 188902 55690
rect 188902 55638 188954 55690
rect 188954 55638 188956 55690
rect 188900 55636 188956 55638
rect 189004 55690 189060 55692
rect 189004 55638 189006 55690
rect 189006 55638 189058 55690
rect 189058 55638 189060 55690
rect 189004 55636 189060 55638
rect 189456 54906 189512 54908
rect 189456 54854 189458 54906
rect 189458 54854 189510 54906
rect 189510 54854 189512 54906
rect 189456 54852 189512 54854
rect 189560 54906 189616 54908
rect 189560 54854 189562 54906
rect 189562 54854 189614 54906
rect 189614 54854 189616 54906
rect 189560 54852 189616 54854
rect 189664 54906 189720 54908
rect 189664 54854 189666 54906
rect 189666 54854 189718 54906
rect 189718 54854 189720 54906
rect 189664 54852 189720 54854
rect 188796 54122 188852 54124
rect 188796 54070 188798 54122
rect 188798 54070 188850 54122
rect 188850 54070 188852 54122
rect 188796 54068 188852 54070
rect 188900 54122 188956 54124
rect 188900 54070 188902 54122
rect 188902 54070 188954 54122
rect 188954 54070 188956 54122
rect 188900 54068 188956 54070
rect 189004 54122 189060 54124
rect 189004 54070 189006 54122
rect 189006 54070 189058 54122
rect 189058 54070 189060 54122
rect 189004 54068 189060 54070
rect 189456 53338 189512 53340
rect 189456 53286 189458 53338
rect 189458 53286 189510 53338
rect 189510 53286 189512 53338
rect 189456 53284 189512 53286
rect 189560 53338 189616 53340
rect 189560 53286 189562 53338
rect 189562 53286 189614 53338
rect 189614 53286 189616 53338
rect 189560 53284 189616 53286
rect 189664 53338 189720 53340
rect 189664 53286 189666 53338
rect 189666 53286 189718 53338
rect 189718 53286 189720 53338
rect 189664 53284 189720 53286
rect 188796 52554 188852 52556
rect 188796 52502 188798 52554
rect 188798 52502 188850 52554
rect 188850 52502 188852 52554
rect 188796 52500 188852 52502
rect 188900 52554 188956 52556
rect 188900 52502 188902 52554
rect 188902 52502 188954 52554
rect 188954 52502 188956 52554
rect 188900 52500 188956 52502
rect 189004 52554 189060 52556
rect 189004 52502 189006 52554
rect 189006 52502 189058 52554
rect 189058 52502 189060 52554
rect 189004 52500 189060 52502
rect 189456 51770 189512 51772
rect 189456 51718 189458 51770
rect 189458 51718 189510 51770
rect 189510 51718 189512 51770
rect 189456 51716 189512 51718
rect 189560 51770 189616 51772
rect 189560 51718 189562 51770
rect 189562 51718 189614 51770
rect 189614 51718 189616 51770
rect 189560 51716 189616 51718
rect 189664 51770 189720 51772
rect 189664 51718 189666 51770
rect 189666 51718 189718 51770
rect 189718 51718 189720 51770
rect 189664 51716 189720 51718
rect 188796 50986 188852 50988
rect 188796 50934 188798 50986
rect 188798 50934 188850 50986
rect 188850 50934 188852 50986
rect 188796 50932 188852 50934
rect 188900 50986 188956 50988
rect 188900 50934 188902 50986
rect 188902 50934 188954 50986
rect 188954 50934 188956 50986
rect 188900 50932 188956 50934
rect 189004 50986 189060 50988
rect 189004 50934 189006 50986
rect 189006 50934 189058 50986
rect 189058 50934 189060 50986
rect 189004 50932 189060 50934
rect 189456 50202 189512 50204
rect 189456 50150 189458 50202
rect 189458 50150 189510 50202
rect 189510 50150 189512 50202
rect 189456 50148 189512 50150
rect 189560 50202 189616 50204
rect 189560 50150 189562 50202
rect 189562 50150 189614 50202
rect 189614 50150 189616 50202
rect 189560 50148 189616 50150
rect 189664 50202 189720 50204
rect 189664 50150 189666 50202
rect 189666 50150 189718 50202
rect 189718 50150 189720 50202
rect 189664 50148 189720 50150
rect 188796 49418 188852 49420
rect 188796 49366 188798 49418
rect 188798 49366 188850 49418
rect 188850 49366 188852 49418
rect 188796 49364 188852 49366
rect 188900 49418 188956 49420
rect 188900 49366 188902 49418
rect 188902 49366 188954 49418
rect 188954 49366 188956 49418
rect 188900 49364 188956 49366
rect 189004 49418 189060 49420
rect 189004 49366 189006 49418
rect 189006 49366 189058 49418
rect 189058 49366 189060 49418
rect 189004 49364 189060 49366
rect 189456 48634 189512 48636
rect 189456 48582 189458 48634
rect 189458 48582 189510 48634
rect 189510 48582 189512 48634
rect 189456 48580 189512 48582
rect 189560 48634 189616 48636
rect 189560 48582 189562 48634
rect 189562 48582 189614 48634
rect 189614 48582 189616 48634
rect 189560 48580 189616 48582
rect 189664 48634 189720 48636
rect 189664 48582 189666 48634
rect 189666 48582 189718 48634
rect 189718 48582 189720 48634
rect 189664 48580 189720 48582
rect 188796 47850 188852 47852
rect 188796 47798 188798 47850
rect 188798 47798 188850 47850
rect 188850 47798 188852 47850
rect 188796 47796 188852 47798
rect 188900 47850 188956 47852
rect 188900 47798 188902 47850
rect 188902 47798 188954 47850
rect 188954 47798 188956 47850
rect 188900 47796 188956 47798
rect 189004 47850 189060 47852
rect 189004 47798 189006 47850
rect 189006 47798 189058 47850
rect 189058 47798 189060 47850
rect 189004 47796 189060 47798
rect 189456 47066 189512 47068
rect 189456 47014 189458 47066
rect 189458 47014 189510 47066
rect 189510 47014 189512 47066
rect 189456 47012 189512 47014
rect 189560 47066 189616 47068
rect 189560 47014 189562 47066
rect 189562 47014 189614 47066
rect 189614 47014 189616 47066
rect 189560 47012 189616 47014
rect 189664 47066 189720 47068
rect 189664 47014 189666 47066
rect 189666 47014 189718 47066
rect 189718 47014 189720 47066
rect 189664 47012 189720 47014
rect 188796 46282 188852 46284
rect 188796 46230 188798 46282
rect 188798 46230 188850 46282
rect 188850 46230 188852 46282
rect 188796 46228 188852 46230
rect 188900 46282 188956 46284
rect 188900 46230 188902 46282
rect 188902 46230 188954 46282
rect 188954 46230 188956 46282
rect 188900 46228 188956 46230
rect 189004 46282 189060 46284
rect 189004 46230 189006 46282
rect 189006 46230 189058 46282
rect 189058 46230 189060 46282
rect 189004 46228 189060 46230
rect 189456 45498 189512 45500
rect 189456 45446 189458 45498
rect 189458 45446 189510 45498
rect 189510 45446 189512 45498
rect 189456 45444 189512 45446
rect 189560 45498 189616 45500
rect 189560 45446 189562 45498
rect 189562 45446 189614 45498
rect 189614 45446 189616 45498
rect 189560 45444 189616 45446
rect 189664 45498 189720 45500
rect 189664 45446 189666 45498
rect 189666 45446 189718 45498
rect 189718 45446 189720 45498
rect 189664 45444 189720 45446
rect 188796 44714 188852 44716
rect 188796 44662 188798 44714
rect 188798 44662 188850 44714
rect 188850 44662 188852 44714
rect 188796 44660 188852 44662
rect 188900 44714 188956 44716
rect 188900 44662 188902 44714
rect 188902 44662 188954 44714
rect 188954 44662 188956 44714
rect 188900 44660 188956 44662
rect 189004 44714 189060 44716
rect 189004 44662 189006 44714
rect 189006 44662 189058 44714
rect 189058 44662 189060 44714
rect 189004 44660 189060 44662
rect 189456 43930 189512 43932
rect 189456 43878 189458 43930
rect 189458 43878 189510 43930
rect 189510 43878 189512 43930
rect 189456 43876 189512 43878
rect 189560 43930 189616 43932
rect 189560 43878 189562 43930
rect 189562 43878 189614 43930
rect 189614 43878 189616 43930
rect 189560 43876 189616 43878
rect 189664 43930 189720 43932
rect 189664 43878 189666 43930
rect 189666 43878 189718 43930
rect 189718 43878 189720 43930
rect 189664 43876 189720 43878
rect 188796 43146 188852 43148
rect 188796 43094 188798 43146
rect 188798 43094 188850 43146
rect 188850 43094 188852 43146
rect 188796 43092 188852 43094
rect 188900 43146 188956 43148
rect 188900 43094 188902 43146
rect 188902 43094 188954 43146
rect 188954 43094 188956 43146
rect 188900 43092 188956 43094
rect 189004 43146 189060 43148
rect 189004 43094 189006 43146
rect 189006 43094 189058 43146
rect 189058 43094 189060 43146
rect 189004 43092 189060 43094
rect 189456 42362 189512 42364
rect 189456 42310 189458 42362
rect 189458 42310 189510 42362
rect 189510 42310 189512 42362
rect 189456 42308 189512 42310
rect 189560 42362 189616 42364
rect 189560 42310 189562 42362
rect 189562 42310 189614 42362
rect 189614 42310 189616 42362
rect 189560 42308 189616 42310
rect 189664 42362 189720 42364
rect 189664 42310 189666 42362
rect 189666 42310 189718 42362
rect 189718 42310 189720 42362
rect 189664 42308 189720 42310
rect 188796 41578 188852 41580
rect 188796 41526 188798 41578
rect 188798 41526 188850 41578
rect 188850 41526 188852 41578
rect 188796 41524 188852 41526
rect 188900 41578 188956 41580
rect 188900 41526 188902 41578
rect 188902 41526 188954 41578
rect 188954 41526 188956 41578
rect 188900 41524 188956 41526
rect 189004 41578 189060 41580
rect 189004 41526 189006 41578
rect 189006 41526 189058 41578
rect 189058 41526 189060 41578
rect 189004 41524 189060 41526
rect 189456 40794 189512 40796
rect 189456 40742 189458 40794
rect 189458 40742 189510 40794
rect 189510 40742 189512 40794
rect 189456 40740 189512 40742
rect 189560 40794 189616 40796
rect 189560 40742 189562 40794
rect 189562 40742 189614 40794
rect 189614 40742 189616 40794
rect 189560 40740 189616 40742
rect 189664 40794 189720 40796
rect 189664 40742 189666 40794
rect 189666 40742 189718 40794
rect 189718 40742 189720 40794
rect 189664 40740 189720 40742
rect 188796 40010 188852 40012
rect 188796 39958 188798 40010
rect 188798 39958 188850 40010
rect 188850 39958 188852 40010
rect 188796 39956 188852 39958
rect 188900 40010 188956 40012
rect 188900 39958 188902 40010
rect 188902 39958 188954 40010
rect 188954 39958 188956 40010
rect 188900 39956 188956 39958
rect 189004 40010 189060 40012
rect 189004 39958 189006 40010
rect 189006 39958 189058 40010
rect 189058 39958 189060 40010
rect 189004 39956 189060 39958
rect 189456 39226 189512 39228
rect 189456 39174 189458 39226
rect 189458 39174 189510 39226
rect 189510 39174 189512 39226
rect 189456 39172 189512 39174
rect 189560 39226 189616 39228
rect 189560 39174 189562 39226
rect 189562 39174 189614 39226
rect 189614 39174 189616 39226
rect 189560 39172 189616 39174
rect 189664 39226 189720 39228
rect 189664 39174 189666 39226
rect 189666 39174 189718 39226
rect 189718 39174 189720 39226
rect 189664 39172 189720 39174
rect 188748 38722 188804 38724
rect 188748 38670 188750 38722
rect 188750 38670 188802 38722
rect 188802 38670 188804 38722
rect 188748 38668 188804 38670
rect 188796 38442 188852 38444
rect 188796 38390 188798 38442
rect 188798 38390 188850 38442
rect 188850 38390 188852 38442
rect 188796 38388 188852 38390
rect 188900 38442 188956 38444
rect 188900 38390 188902 38442
rect 188902 38390 188954 38442
rect 188954 38390 188956 38442
rect 188900 38388 188956 38390
rect 189004 38442 189060 38444
rect 189004 38390 189006 38442
rect 189006 38390 189058 38442
rect 189058 38390 189060 38442
rect 189004 38388 189060 38390
rect 189456 37658 189512 37660
rect 189456 37606 189458 37658
rect 189458 37606 189510 37658
rect 189510 37606 189512 37658
rect 189456 37604 189512 37606
rect 189560 37658 189616 37660
rect 189560 37606 189562 37658
rect 189562 37606 189614 37658
rect 189614 37606 189616 37658
rect 189560 37604 189616 37606
rect 189664 37658 189720 37660
rect 189664 37606 189666 37658
rect 189666 37606 189718 37658
rect 189718 37606 189720 37658
rect 189664 37604 189720 37606
rect 188796 36874 188852 36876
rect 188796 36822 188798 36874
rect 188798 36822 188850 36874
rect 188850 36822 188852 36874
rect 188796 36820 188852 36822
rect 188900 36874 188956 36876
rect 188900 36822 188902 36874
rect 188902 36822 188954 36874
rect 188954 36822 188956 36874
rect 188900 36820 188956 36822
rect 189004 36874 189060 36876
rect 189004 36822 189006 36874
rect 189006 36822 189058 36874
rect 189058 36822 189060 36874
rect 189004 36820 189060 36822
rect 189456 36090 189512 36092
rect 189456 36038 189458 36090
rect 189458 36038 189510 36090
rect 189510 36038 189512 36090
rect 189456 36036 189512 36038
rect 189560 36090 189616 36092
rect 189560 36038 189562 36090
rect 189562 36038 189614 36090
rect 189614 36038 189616 36090
rect 189560 36036 189616 36038
rect 189664 36090 189720 36092
rect 189664 36038 189666 36090
rect 189666 36038 189718 36090
rect 189718 36038 189720 36090
rect 189664 36036 189720 36038
rect 188796 35306 188852 35308
rect 188796 35254 188798 35306
rect 188798 35254 188850 35306
rect 188850 35254 188852 35306
rect 188796 35252 188852 35254
rect 188900 35306 188956 35308
rect 188900 35254 188902 35306
rect 188902 35254 188954 35306
rect 188954 35254 188956 35306
rect 188900 35252 188956 35254
rect 189004 35306 189060 35308
rect 189004 35254 189006 35306
rect 189006 35254 189058 35306
rect 189058 35254 189060 35306
rect 189004 35252 189060 35254
rect 189456 34522 189512 34524
rect 189456 34470 189458 34522
rect 189458 34470 189510 34522
rect 189510 34470 189512 34522
rect 189456 34468 189512 34470
rect 189560 34522 189616 34524
rect 189560 34470 189562 34522
rect 189562 34470 189614 34522
rect 189614 34470 189616 34522
rect 189560 34468 189616 34470
rect 189664 34522 189720 34524
rect 189664 34470 189666 34522
rect 189666 34470 189718 34522
rect 189718 34470 189720 34522
rect 189664 34468 189720 34470
rect 188796 33738 188852 33740
rect 188796 33686 188798 33738
rect 188798 33686 188850 33738
rect 188850 33686 188852 33738
rect 188796 33684 188852 33686
rect 188900 33738 188956 33740
rect 188900 33686 188902 33738
rect 188902 33686 188954 33738
rect 188954 33686 188956 33738
rect 188900 33684 188956 33686
rect 189004 33738 189060 33740
rect 189004 33686 189006 33738
rect 189006 33686 189058 33738
rect 189058 33686 189060 33738
rect 189004 33684 189060 33686
rect 189456 32954 189512 32956
rect 189456 32902 189458 32954
rect 189458 32902 189510 32954
rect 189510 32902 189512 32954
rect 189456 32900 189512 32902
rect 189560 32954 189616 32956
rect 189560 32902 189562 32954
rect 189562 32902 189614 32954
rect 189614 32902 189616 32954
rect 189560 32900 189616 32902
rect 189664 32954 189720 32956
rect 189664 32902 189666 32954
rect 189666 32902 189718 32954
rect 189718 32902 189720 32954
rect 189664 32900 189720 32902
rect 188796 32170 188852 32172
rect 188796 32118 188798 32170
rect 188798 32118 188850 32170
rect 188850 32118 188852 32170
rect 188796 32116 188852 32118
rect 188900 32170 188956 32172
rect 188900 32118 188902 32170
rect 188902 32118 188954 32170
rect 188954 32118 188956 32170
rect 188900 32116 188956 32118
rect 189004 32170 189060 32172
rect 189004 32118 189006 32170
rect 189006 32118 189058 32170
rect 189058 32118 189060 32170
rect 189004 32116 189060 32118
rect 189456 31386 189512 31388
rect 189456 31334 189458 31386
rect 189458 31334 189510 31386
rect 189510 31334 189512 31386
rect 189456 31332 189512 31334
rect 189560 31386 189616 31388
rect 189560 31334 189562 31386
rect 189562 31334 189614 31386
rect 189614 31334 189616 31386
rect 189560 31332 189616 31334
rect 189664 31386 189720 31388
rect 189664 31334 189666 31386
rect 189666 31334 189718 31386
rect 189718 31334 189720 31386
rect 189664 31332 189720 31334
rect 188796 30602 188852 30604
rect 188796 30550 188798 30602
rect 188798 30550 188850 30602
rect 188850 30550 188852 30602
rect 188796 30548 188852 30550
rect 188900 30602 188956 30604
rect 188900 30550 188902 30602
rect 188902 30550 188954 30602
rect 188954 30550 188956 30602
rect 188900 30548 188956 30550
rect 189004 30602 189060 30604
rect 189004 30550 189006 30602
rect 189006 30550 189058 30602
rect 189058 30550 189060 30602
rect 189004 30548 189060 30550
rect 189456 29818 189512 29820
rect 189456 29766 189458 29818
rect 189458 29766 189510 29818
rect 189510 29766 189512 29818
rect 189456 29764 189512 29766
rect 189560 29818 189616 29820
rect 189560 29766 189562 29818
rect 189562 29766 189614 29818
rect 189614 29766 189616 29818
rect 189560 29764 189616 29766
rect 189664 29818 189720 29820
rect 189664 29766 189666 29818
rect 189666 29766 189718 29818
rect 189718 29766 189720 29818
rect 189664 29764 189720 29766
rect 188796 29034 188852 29036
rect 188796 28982 188798 29034
rect 188798 28982 188850 29034
rect 188850 28982 188852 29034
rect 188796 28980 188852 28982
rect 188900 29034 188956 29036
rect 188900 28982 188902 29034
rect 188902 28982 188954 29034
rect 188954 28982 188956 29034
rect 188900 28980 188956 28982
rect 189004 29034 189060 29036
rect 189004 28982 189006 29034
rect 189006 28982 189058 29034
rect 189058 28982 189060 29034
rect 189004 28980 189060 28982
rect 189456 28250 189512 28252
rect 189456 28198 189458 28250
rect 189458 28198 189510 28250
rect 189510 28198 189512 28250
rect 189456 28196 189512 28198
rect 189560 28250 189616 28252
rect 189560 28198 189562 28250
rect 189562 28198 189614 28250
rect 189614 28198 189616 28250
rect 189560 28196 189616 28198
rect 189664 28250 189720 28252
rect 189664 28198 189666 28250
rect 189666 28198 189718 28250
rect 189718 28198 189720 28250
rect 189664 28196 189720 28198
rect 188796 27466 188852 27468
rect 188796 27414 188798 27466
rect 188798 27414 188850 27466
rect 188850 27414 188852 27466
rect 188796 27412 188852 27414
rect 188900 27466 188956 27468
rect 188900 27414 188902 27466
rect 188902 27414 188954 27466
rect 188954 27414 188956 27466
rect 188900 27412 188956 27414
rect 189004 27466 189060 27468
rect 189004 27414 189006 27466
rect 189006 27414 189058 27466
rect 189058 27414 189060 27466
rect 189004 27412 189060 27414
rect 189456 26682 189512 26684
rect 189456 26630 189458 26682
rect 189458 26630 189510 26682
rect 189510 26630 189512 26682
rect 189456 26628 189512 26630
rect 189560 26682 189616 26684
rect 189560 26630 189562 26682
rect 189562 26630 189614 26682
rect 189614 26630 189616 26682
rect 189560 26628 189616 26630
rect 189664 26682 189720 26684
rect 189664 26630 189666 26682
rect 189666 26630 189718 26682
rect 189718 26630 189720 26682
rect 189664 26628 189720 26630
rect 188796 25898 188852 25900
rect 188796 25846 188798 25898
rect 188798 25846 188850 25898
rect 188850 25846 188852 25898
rect 188796 25844 188852 25846
rect 188900 25898 188956 25900
rect 188900 25846 188902 25898
rect 188902 25846 188954 25898
rect 188954 25846 188956 25898
rect 188900 25844 188956 25846
rect 189004 25898 189060 25900
rect 189004 25846 189006 25898
rect 189006 25846 189058 25898
rect 189058 25846 189060 25898
rect 189004 25844 189060 25846
rect 187292 25564 187348 25620
rect 204316 154140 204372 154196
rect 196588 29372 196644 29428
rect 201068 146242 201124 146244
rect 201068 146190 201070 146242
rect 201070 146190 201122 146242
rect 201122 146190 201124 146242
rect 201068 146188 201124 146190
rect 201740 146242 201796 146244
rect 201740 146190 201742 146242
rect 201742 146190 201794 146242
rect 201794 146190 201796 146242
rect 201740 146188 201796 146190
rect 204092 145404 204148 145460
rect 203756 127932 203812 127988
rect 204092 119308 204148 119364
rect 202188 118636 202244 118692
rect 203756 118690 203812 118692
rect 203756 118638 203758 118690
rect 203758 118638 203810 118690
rect 203810 118638 203812 118690
rect 203756 118636 203812 118638
rect 201180 93714 201236 93716
rect 201180 93662 201182 93714
rect 201182 93662 201234 93714
rect 201234 93662 201236 93714
rect 201180 93660 201236 93662
rect 201180 67058 201236 67060
rect 201180 67006 201182 67058
rect 201182 67006 201234 67058
rect 201234 67006 201236 67058
rect 201180 67004 201236 67006
rect 201404 40962 201460 40964
rect 201404 40910 201406 40962
rect 201406 40910 201458 40962
rect 201458 40910 201460 40962
rect 201404 40908 201460 40910
rect 201068 27804 201124 27860
rect 204316 101724 204372 101780
rect 203980 93660 204036 93716
rect 203196 92988 203252 93044
rect 204316 75570 204372 75572
rect 204316 75518 204318 75570
rect 204318 75518 204370 75570
rect 204370 75518 204372 75570
rect 204316 75516 204372 75518
rect 203980 67004 204036 67060
rect 203196 66780 203252 66836
rect 203756 49308 203812 49364
rect 204092 40572 204148 40628
rect 202412 27692 202468 27748
rect 190652 25340 190708 25396
rect 189456 25114 189512 25116
rect 189456 25062 189458 25114
rect 189458 25062 189510 25114
rect 189510 25062 189512 25114
rect 189456 25060 189512 25062
rect 189560 25114 189616 25116
rect 189560 25062 189562 25114
rect 189562 25062 189614 25114
rect 189614 25062 189616 25114
rect 189560 25060 189616 25062
rect 189664 25114 189720 25116
rect 189664 25062 189666 25114
rect 189666 25062 189718 25114
rect 189718 25062 189720 25114
rect 189664 25060 189720 25062
rect 188796 24330 188852 24332
rect 188796 24278 188798 24330
rect 188798 24278 188850 24330
rect 188850 24278 188852 24330
rect 188796 24276 188852 24278
rect 188900 24330 188956 24332
rect 188900 24278 188902 24330
rect 188902 24278 188954 24330
rect 188954 24278 188956 24330
rect 188900 24276 188956 24278
rect 189004 24330 189060 24332
rect 189004 24278 189006 24330
rect 189006 24278 189058 24330
rect 189058 24278 189060 24330
rect 189004 24276 189060 24278
rect 189456 23546 189512 23548
rect 189456 23494 189458 23546
rect 189458 23494 189510 23546
rect 189510 23494 189512 23546
rect 189456 23492 189512 23494
rect 189560 23546 189616 23548
rect 189560 23494 189562 23546
rect 189562 23494 189614 23546
rect 189614 23494 189616 23546
rect 189560 23492 189616 23494
rect 189664 23546 189720 23548
rect 189664 23494 189666 23546
rect 189666 23494 189718 23546
rect 189718 23494 189720 23546
rect 189664 23492 189720 23494
rect 204316 23100 204372 23156
rect 188796 22762 188852 22764
rect 188796 22710 188798 22762
rect 188798 22710 188850 22762
rect 188850 22710 188852 22762
rect 188796 22708 188852 22710
rect 188900 22762 188956 22764
rect 188900 22710 188902 22762
rect 188902 22710 188954 22762
rect 188954 22710 188956 22762
rect 188900 22708 188956 22710
rect 189004 22762 189060 22764
rect 189004 22710 189006 22762
rect 189006 22710 189058 22762
rect 189058 22710 189060 22762
rect 189004 22708 189060 22710
rect 189456 21978 189512 21980
rect 189456 21926 189458 21978
rect 189458 21926 189510 21978
rect 189510 21926 189512 21978
rect 189456 21924 189512 21926
rect 189560 21978 189616 21980
rect 189560 21926 189562 21978
rect 189562 21926 189614 21978
rect 189614 21926 189616 21978
rect 189560 21924 189616 21926
rect 189664 21978 189720 21980
rect 189664 21926 189666 21978
rect 189666 21926 189718 21978
rect 189718 21926 189720 21978
rect 189664 21924 189720 21926
rect 188796 21194 188852 21196
rect 188796 21142 188798 21194
rect 188798 21142 188850 21194
rect 188850 21142 188852 21194
rect 188796 21140 188852 21142
rect 188900 21194 188956 21196
rect 188900 21142 188902 21194
rect 188902 21142 188954 21194
rect 188954 21142 188956 21194
rect 188900 21140 188956 21142
rect 189004 21194 189060 21196
rect 189004 21142 189006 21194
rect 189006 21142 189058 21194
rect 189058 21142 189060 21194
rect 189004 21140 189060 21142
rect 154588 20412 154644 20468
rect 189456 20410 189512 20412
rect 189456 20358 189458 20410
rect 189458 20358 189510 20410
rect 189510 20358 189512 20410
rect 189456 20356 189512 20358
rect 189560 20410 189616 20412
rect 189560 20358 189562 20410
rect 189562 20358 189614 20410
rect 189614 20358 189616 20410
rect 189560 20356 189616 20358
rect 189664 20410 189720 20412
rect 189664 20358 189666 20410
rect 189666 20358 189718 20410
rect 189718 20358 189720 20410
rect 189664 20356 189720 20358
rect 188796 19626 188852 19628
rect 188796 19574 188798 19626
rect 188798 19574 188850 19626
rect 188850 19574 188852 19626
rect 188796 19572 188852 19574
rect 188900 19626 188956 19628
rect 188900 19574 188902 19626
rect 188902 19574 188954 19626
rect 188954 19574 188956 19626
rect 188900 19572 188956 19574
rect 189004 19626 189060 19628
rect 189004 19574 189006 19626
rect 189006 19574 189058 19626
rect 189058 19574 189060 19626
rect 189004 19572 189060 19574
rect 189456 18842 189512 18844
rect 189456 18790 189458 18842
rect 189458 18790 189510 18842
rect 189510 18790 189512 18842
rect 189456 18788 189512 18790
rect 189560 18842 189616 18844
rect 189560 18790 189562 18842
rect 189562 18790 189614 18842
rect 189614 18790 189616 18842
rect 189560 18788 189616 18790
rect 189664 18842 189720 18844
rect 189664 18790 189666 18842
rect 189666 18790 189718 18842
rect 189718 18790 189720 18842
rect 189664 18788 189720 18790
rect 188796 18058 188852 18060
rect 188796 18006 188798 18058
rect 188798 18006 188850 18058
rect 188850 18006 188852 18058
rect 188796 18004 188852 18006
rect 188900 18058 188956 18060
rect 188900 18006 188902 18058
rect 188902 18006 188954 18058
rect 188954 18006 188956 18058
rect 188900 18004 188956 18006
rect 189004 18058 189060 18060
rect 189004 18006 189006 18058
rect 189006 18006 189058 18058
rect 189058 18006 189060 18058
rect 189004 18004 189060 18006
rect 158736 17274 158792 17276
rect 158736 17222 158738 17274
rect 158738 17222 158790 17274
rect 158790 17222 158792 17274
rect 158736 17220 158792 17222
rect 158840 17274 158896 17276
rect 158840 17222 158842 17274
rect 158842 17222 158894 17274
rect 158894 17222 158896 17274
rect 158840 17220 158896 17222
rect 158944 17274 159000 17276
rect 158944 17222 158946 17274
rect 158946 17222 158998 17274
rect 158998 17222 159000 17274
rect 158944 17220 159000 17222
rect 189456 17274 189512 17276
rect 189456 17222 189458 17274
rect 189458 17222 189510 17274
rect 189510 17222 189512 17274
rect 189456 17220 189512 17222
rect 189560 17274 189616 17276
rect 189560 17222 189562 17274
rect 189562 17222 189614 17274
rect 189614 17222 189616 17274
rect 189560 17220 189616 17222
rect 189664 17274 189720 17276
rect 189664 17222 189666 17274
rect 189666 17222 189718 17274
rect 189718 17222 189720 17274
rect 189664 17220 189720 17222
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 35856 15706 35912 15708
rect 35856 15654 35858 15706
rect 35858 15654 35910 15706
rect 35910 15654 35912 15706
rect 35856 15652 35912 15654
rect 35960 15706 36016 15708
rect 35960 15654 35962 15706
rect 35962 15654 36014 15706
rect 36014 15654 36016 15706
rect 35960 15652 36016 15654
rect 36064 15706 36120 15708
rect 36064 15654 36066 15706
rect 36066 15654 36118 15706
rect 36118 15654 36120 15706
rect 36064 15652 36120 15654
rect 66576 15706 66632 15708
rect 66576 15654 66578 15706
rect 66578 15654 66630 15706
rect 66630 15654 66632 15706
rect 66576 15652 66632 15654
rect 66680 15706 66736 15708
rect 66680 15654 66682 15706
rect 66682 15654 66734 15706
rect 66734 15654 66736 15706
rect 66680 15652 66736 15654
rect 66784 15706 66840 15708
rect 66784 15654 66786 15706
rect 66786 15654 66838 15706
rect 66838 15654 66840 15706
rect 66784 15652 66840 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 125580 16882 125636 16884
rect 125580 16830 125582 16882
rect 125582 16830 125634 16882
rect 125634 16830 125636 16882
rect 125580 16828 125636 16830
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 127356 16490 127412 16492
rect 127356 16438 127358 16490
rect 127358 16438 127410 16490
rect 127410 16438 127412 16490
rect 127356 16436 127412 16438
rect 127460 16490 127516 16492
rect 127460 16438 127462 16490
rect 127462 16438 127514 16490
rect 127514 16438 127516 16490
rect 127460 16436 127516 16438
rect 127564 16490 127620 16492
rect 127564 16438 127566 16490
rect 127566 16438 127618 16490
rect 127618 16438 127620 16490
rect 127564 16436 127620 16438
rect 158076 16490 158132 16492
rect 158076 16438 158078 16490
rect 158078 16438 158130 16490
rect 158130 16438 158132 16490
rect 158076 16436 158132 16438
rect 158180 16490 158236 16492
rect 158180 16438 158182 16490
rect 158182 16438 158234 16490
rect 158234 16438 158236 16490
rect 158180 16436 158236 16438
rect 158284 16490 158340 16492
rect 158284 16438 158286 16490
rect 158286 16438 158338 16490
rect 158338 16438 158340 16490
rect 158284 16436 158340 16438
rect 188796 16490 188852 16492
rect 188796 16438 188798 16490
rect 188798 16438 188850 16490
rect 188850 16438 188852 16490
rect 188796 16436 188852 16438
rect 188900 16490 188956 16492
rect 188900 16438 188902 16490
rect 188902 16438 188954 16490
rect 188954 16438 188956 16490
rect 188900 16436 188956 16438
rect 189004 16490 189060 16492
rect 189004 16438 189006 16490
rect 189006 16438 189058 16490
rect 189058 16438 189060 16490
rect 189004 16436 189060 16438
rect 97296 15706 97352 15708
rect 97296 15654 97298 15706
rect 97298 15654 97350 15706
rect 97350 15654 97352 15706
rect 97296 15652 97352 15654
rect 97400 15706 97456 15708
rect 97400 15654 97402 15706
rect 97402 15654 97454 15706
rect 97454 15654 97456 15706
rect 97400 15652 97456 15654
rect 97504 15706 97560 15708
rect 97504 15654 97506 15706
rect 97506 15654 97558 15706
rect 97558 15654 97560 15706
rect 97504 15652 97560 15654
rect 128016 15706 128072 15708
rect 128016 15654 128018 15706
rect 128018 15654 128070 15706
rect 128070 15654 128072 15706
rect 128016 15652 128072 15654
rect 128120 15706 128176 15708
rect 128120 15654 128122 15706
rect 128122 15654 128174 15706
rect 128174 15654 128176 15706
rect 128120 15652 128176 15654
rect 128224 15706 128280 15708
rect 128224 15654 128226 15706
rect 128226 15654 128278 15706
rect 128278 15654 128280 15706
rect 128224 15652 128280 15654
rect 158736 15706 158792 15708
rect 158736 15654 158738 15706
rect 158738 15654 158790 15706
rect 158790 15654 158792 15706
rect 158736 15652 158792 15654
rect 158840 15706 158896 15708
rect 158840 15654 158842 15706
rect 158842 15654 158894 15706
rect 158894 15654 158896 15706
rect 158840 15652 158896 15654
rect 158944 15706 159000 15708
rect 158944 15654 158946 15706
rect 158946 15654 158998 15706
rect 158998 15654 159000 15706
rect 158944 15652 159000 15654
rect 189456 15706 189512 15708
rect 189456 15654 189458 15706
rect 189458 15654 189510 15706
rect 189510 15654 189512 15706
rect 189456 15652 189512 15654
rect 189560 15706 189616 15708
rect 189560 15654 189562 15706
rect 189562 15654 189614 15706
rect 189614 15654 189616 15706
rect 189560 15652 189616 15654
rect 189664 15706 189720 15708
rect 189664 15654 189666 15706
rect 189666 15654 189718 15706
rect 189718 15654 189720 15706
rect 189664 15652 189720 15654
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 127356 14922 127412 14924
rect 127356 14870 127358 14922
rect 127358 14870 127410 14922
rect 127410 14870 127412 14922
rect 127356 14868 127412 14870
rect 127460 14922 127516 14924
rect 127460 14870 127462 14922
rect 127462 14870 127514 14922
rect 127514 14870 127516 14922
rect 127460 14868 127516 14870
rect 127564 14922 127620 14924
rect 127564 14870 127566 14922
rect 127566 14870 127618 14922
rect 127618 14870 127620 14922
rect 127564 14868 127620 14870
rect 158076 14922 158132 14924
rect 158076 14870 158078 14922
rect 158078 14870 158130 14922
rect 158130 14870 158132 14922
rect 158076 14868 158132 14870
rect 158180 14922 158236 14924
rect 158180 14870 158182 14922
rect 158182 14870 158234 14922
rect 158234 14870 158236 14922
rect 158180 14868 158236 14870
rect 158284 14922 158340 14924
rect 158284 14870 158286 14922
rect 158286 14870 158338 14922
rect 158338 14870 158340 14922
rect 158284 14868 158340 14870
rect 188796 14922 188852 14924
rect 188796 14870 188798 14922
rect 188798 14870 188850 14922
rect 188850 14870 188852 14922
rect 188796 14868 188852 14870
rect 188900 14922 188956 14924
rect 188900 14870 188902 14922
rect 188902 14870 188954 14922
rect 188954 14870 188956 14922
rect 188900 14868 188956 14870
rect 189004 14922 189060 14924
rect 189004 14870 189006 14922
rect 189006 14870 189058 14922
rect 189058 14870 189060 14922
rect 189004 14868 189060 14870
rect 67900 14476 67956 14532
rect 201740 14530 201796 14532
rect 201740 14478 201742 14530
rect 201742 14478 201794 14530
rect 201794 14478 201796 14530
rect 201740 14476 201796 14478
rect 204092 14364 204148 14420
rect 204316 14476 204372 14532
rect 35856 14138 35912 14140
rect 35856 14086 35858 14138
rect 35858 14086 35910 14138
rect 35910 14086 35912 14138
rect 35856 14084 35912 14086
rect 35960 14138 36016 14140
rect 35960 14086 35962 14138
rect 35962 14086 36014 14138
rect 36014 14086 36016 14138
rect 35960 14084 36016 14086
rect 36064 14138 36120 14140
rect 36064 14086 36066 14138
rect 36066 14086 36118 14138
rect 36118 14086 36120 14138
rect 36064 14084 36120 14086
rect 66576 14138 66632 14140
rect 66576 14086 66578 14138
rect 66578 14086 66630 14138
rect 66630 14086 66632 14138
rect 66576 14084 66632 14086
rect 66680 14138 66736 14140
rect 66680 14086 66682 14138
rect 66682 14086 66734 14138
rect 66734 14086 66736 14138
rect 66680 14084 66736 14086
rect 66784 14138 66840 14140
rect 66784 14086 66786 14138
rect 66786 14086 66838 14138
rect 66838 14086 66840 14138
rect 66784 14084 66840 14086
rect 97296 14138 97352 14140
rect 97296 14086 97298 14138
rect 97298 14086 97350 14138
rect 97350 14086 97352 14138
rect 97296 14084 97352 14086
rect 97400 14138 97456 14140
rect 97400 14086 97402 14138
rect 97402 14086 97454 14138
rect 97454 14086 97456 14138
rect 97400 14084 97456 14086
rect 97504 14138 97560 14140
rect 97504 14086 97506 14138
rect 97506 14086 97558 14138
rect 97558 14086 97560 14138
rect 97504 14084 97560 14086
rect 128016 14138 128072 14140
rect 128016 14086 128018 14138
rect 128018 14086 128070 14138
rect 128070 14086 128072 14138
rect 128016 14084 128072 14086
rect 128120 14138 128176 14140
rect 128120 14086 128122 14138
rect 128122 14086 128174 14138
rect 128174 14086 128176 14138
rect 128120 14084 128176 14086
rect 128224 14138 128280 14140
rect 128224 14086 128226 14138
rect 128226 14086 128278 14138
rect 128278 14086 128280 14138
rect 128224 14084 128280 14086
rect 158736 14138 158792 14140
rect 158736 14086 158738 14138
rect 158738 14086 158790 14138
rect 158790 14086 158792 14138
rect 158736 14084 158792 14086
rect 158840 14138 158896 14140
rect 158840 14086 158842 14138
rect 158842 14086 158894 14138
rect 158894 14086 158896 14138
rect 158840 14084 158896 14086
rect 158944 14138 159000 14140
rect 158944 14086 158946 14138
rect 158946 14086 158998 14138
rect 158998 14086 159000 14138
rect 158944 14084 159000 14086
rect 189456 14138 189512 14140
rect 189456 14086 189458 14138
rect 189458 14086 189510 14138
rect 189510 14086 189512 14138
rect 189456 14084 189512 14086
rect 189560 14138 189616 14140
rect 189560 14086 189562 14138
rect 189562 14086 189614 14138
rect 189614 14086 189616 14138
rect 189560 14084 189616 14086
rect 189664 14138 189720 14140
rect 189664 14086 189666 14138
rect 189666 14086 189718 14138
rect 189718 14086 189720 14138
rect 189664 14084 189720 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 127356 13354 127412 13356
rect 127356 13302 127358 13354
rect 127358 13302 127410 13354
rect 127410 13302 127412 13354
rect 127356 13300 127412 13302
rect 127460 13354 127516 13356
rect 127460 13302 127462 13354
rect 127462 13302 127514 13354
rect 127514 13302 127516 13354
rect 127460 13300 127516 13302
rect 127564 13354 127620 13356
rect 127564 13302 127566 13354
rect 127566 13302 127618 13354
rect 127618 13302 127620 13354
rect 127564 13300 127620 13302
rect 158076 13354 158132 13356
rect 158076 13302 158078 13354
rect 158078 13302 158130 13354
rect 158130 13302 158132 13354
rect 158076 13300 158132 13302
rect 158180 13354 158236 13356
rect 158180 13302 158182 13354
rect 158182 13302 158234 13354
rect 158234 13302 158236 13354
rect 158180 13300 158236 13302
rect 158284 13354 158340 13356
rect 158284 13302 158286 13354
rect 158286 13302 158338 13354
rect 158338 13302 158340 13354
rect 158284 13300 158340 13302
rect 188796 13354 188852 13356
rect 188796 13302 188798 13354
rect 188798 13302 188850 13354
rect 188850 13302 188852 13354
rect 188796 13300 188852 13302
rect 188900 13354 188956 13356
rect 188900 13302 188902 13354
rect 188902 13302 188954 13354
rect 188954 13302 188956 13354
rect 188900 13300 188956 13302
rect 189004 13354 189060 13356
rect 189004 13302 189006 13354
rect 189006 13302 189058 13354
rect 189058 13302 189060 13354
rect 189004 13300 189060 13302
rect 35856 12570 35912 12572
rect 35856 12518 35858 12570
rect 35858 12518 35910 12570
rect 35910 12518 35912 12570
rect 35856 12516 35912 12518
rect 35960 12570 36016 12572
rect 35960 12518 35962 12570
rect 35962 12518 36014 12570
rect 36014 12518 36016 12570
rect 35960 12516 36016 12518
rect 36064 12570 36120 12572
rect 36064 12518 36066 12570
rect 36066 12518 36118 12570
rect 36118 12518 36120 12570
rect 36064 12516 36120 12518
rect 66576 12570 66632 12572
rect 66576 12518 66578 12570
rect 66578 12518 66630 12570
rect 66630 12518 66632 12570
rect 66576 12516 66632 12518
rect 66680 12570 66736 12572
rect 66680 12518 66682 12570
rect 66682 12518 66734 12570
rect 66734 12518 66736 12570
rect 66680 12516 66736 12518
rect 66784 12570 66840 12572
rect 66784 12518 66786 12570
rect 66786 12518 66838 12570
rect 66838 12518 66840 12570
rect 66784 12516 66840 12518
rect 97296 12570 97352 12572
rect 97296 12518 97298 12570
rect 97298 12518 97350 12570
rect 97350 12518 97352 12570
rect 97296 12516 97352 12518
rect 97400 12570 97456 12572
rect 97400 12518 97402 12570
rect 97402 12518 97454 12570
rect 97454 12518 97456 12570
rect 97400 12516 97456 12518
rect 97504 12570 97560 12572
rect 97504 12518 97506 12570
rect 97506 12518 97558 12570
rect 97558 12518 97560 12570
rect 97504 12516 97560 12518
rect 128016 12570 128072 12572
rect 128016 12518 128018 12570
rect 128018 12518 128070 12570
rect 128070 12518 128072 12570
rect 128016 12516 128072 12518
rect 128120 12570 128176 12572
rect 128120 12518 128122 12570
rect 128122 12518 128174 12570
rect 128174 12518 128176 12570
rect 128120 12516 128176 12518
rect 128224 12570 128280 12572
rect 128224 12518 128226 12570
rect 128226 12518 128278 12570
rect 128278 12518 128280 12570
rect 128224 12516 128280 12518
rect 158736 12570 158792 12572
rect 158736 12518 158738 12570
rect 158738 12518 158790 12570
rect 158790 12518 158792 12570
rect 158736 12516 158792 12518
rect 158840 12570 158896 12572
rect 158840 12518 158842 12570
rect 158842 12518 158894 12570
rect 158894 12518 158896 12570
rect 158840 12516 158896 12518
rect 158944 12570 159000 12572
rect 158944 12518 158946 12570
rect 158946 12518 158998 12570
rect 158998 12518 159000 12570
rect 158944 12516 159000 12518
rect 189456 12570 189512 12572
rect 189456 12518 189458 12570
rect 189458 12518 189510 12570
rect 189510 12518 189512 12570
rect 189456 12516 189512 12518
rect 189560 12570 189616 12572
rect 189560 12518 189562 12570
rect 189562 12518 189614 12570
rect 189614 12518 189616 12570
rect 189560 12516 189616 12518
rect 189664 12570 189720 12572
rect 189664 12518 189666 12570
rect 189666 12518 189718 12570
rect 189718 12518 189720 12570
rect 189664 12516 189720 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 127356 11786 127412 11788
rect 127356 11734 127358 11786
rect 127358 11734 127410 11786
rect 127410 11734 127412 11786
rect 127356 11732 127412 11734
rect 127460 11786 127516 11788
rect 127460 11734 127462 11786
rect 127462 11734 127514 11786
rect 127514 11734 127516 11786
rect 127460 11732 127516 11734
rect 127564 11786 127620 11788
rect 127564 11734 127566 11786
rect 127566 11734 127618 11786
rect 127618 11734 127620 11786
rect 127564 11732 127620 11734
rect 158076 11786 158132 11788
rect 158076 11734 158078 11786
rect 158078 11734 158130 11786
rect 158130 11734 158132 11786
rect 158076 11732 158132 11734
rect 158180 11786 158236 11788
rect 158180 11734 158182 11786
rect 158182 11734 158234 11786
rect 158234 11734 158236 11786
rect 158180 11732 158236 11734
rect 158284 11786 158340 11788
rect 158284 11734 158286 11786
rect 158286 11734 158338 11786
rect 158338 11734 158340 11786
rect 158284 11732 158340 11734
rect 188796 11786 188852 11788
rect 188796 11734 188798 11786
rect 188798 11734 188850 11786
rect 188850 11734 188852 11786
rect 188796 11732 188852 11734
rect 188900 11786 188956 11788
rect 188900 11734 188902 11786
rect 188902 11734 188954 11786
rect 188954 11734 188956 11786
rect 188900 11732 188956 11734
rect 189004 11786 189060 11788
rect 189004 11734 189006 11786
rect 189006 11734 189058 11786
rect 189058 11734 189060 11786
rect 189004 11732 189060 11734
rect 35856 11002 35912 11004
rect 35856 10950 35858 11002
rect 35858 10950 35910 11002
rect 35910 10950 35912 11002
rect 35856 10948 35912 10950
rect 35960 11002 36016 11004
rect 35960 10950 35962 11002
rect 35962 10950 36014 11002
rect 36014 10950 36016 11002
rect 35960 10948 36016 10950
rect 36064 11002 36120 11004
rect 36064 10950 36066 11002
rect 36066 10950 36118 11002
rect 36118 10950 36120 11002
rect 36064 10948 36120 10950
rect 66576 11002 66632 11004
rect 66576 10950 66578 11002
rect 66578 10950 66630 11002
rect 66630 10950 66632 11002
rect 66576 10948 66632 10950
rect 66680 11002 66736 11004
rect 66680 10950 66682 11002
rect 66682 10950 66734 11002
rect 66734 10950 66736 11002
rect 66680 10948 66736 10950
rect 66784 11002 66840 11004
rect 66784 10950 66786 11002
rect 66786 10950 66838 11002
rect 66838 10950 66840 11002
rect 66784 10948 66840 10950
rect 97296 11002 97352 11004
rect 97296 10950 97298 11002
rect 97298 10950 97350 11002
rect 97350 10950 97352 11002
rect 97296 10948 97352 10950
rect 97400 11002 97456 11004
rect 97400 10950 97402 11002
rect 97402 10950 97454 11002
rect 97454 10950 97456 11002
rect 97400 10948 97456 10950
rect 97504 11002 97560 11004
rect 97504 10950 97506 11002
rect 97506 10950 97558 11002
rect 97558 10950 97560 11002
rect 97504 10948 97560 10950
rect 128016 11002 128072 11004
rect 128016 10950 128018 11002
rect 128018 10950 128070 11002
rect 128070 10950 128072 11002
rect 128016 10948 128072 10950
rect 128120 11002 128176 11004
rect 128120 10950 128122 11002
rect 128122 10950 128174 11002
rect 128174 10950 128176 11002
rect 128120 10948 128176 10950
rect 128224 11002 128280 11004
rect 128224 10950 128226 11002
rect 128226 10950 128278 11002
rect 128278 10950 128280 11002
rect 128224 10948 128280 10950
rect 158736 11002 158792 11004
rect 158736 10950 158738 11002
rect 158738 10950 158790 11002
rect 158790 10950 158792 11002
rect 158736 10948 158792 10950
rect 158840 11002 158896 11004
rect 158840 10950 158842 11002
rect 158842 10950 158894 11002
rect 158894 10950 158896 11002
rect 158840 10948 158896 10950
rect 158944 11002 159000 11004
rect 158944 10950 158946 11002
rect 158946 10950 158998 11002
rect 158998 10950 159000 11002
rect 158944 10948 159000 10950
rect 189456 11002 189512 11004
rect 189456 10950 189458 11002
rect 189458 10950 189510 11002
rect 189510 10950 189512 11002
rect 189456 10948 189512 10950
rect 189560 11002 189616 11004
rect 189560 10950 189562 11002
rect 189562 10950 189614 11002
rect 189614 10950 189616 11002
rect 189560 10948 189616 10950
rect 189664 11002 189720 11004
rect 189664 10950 189666 11002
rect 189666 10950 189718 11002
rect 189718 10950 189720 11002
rect 189664 10948 189720 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 127356 10218 127412 10220
rect 127356 10166 127358 10218
rect 127358 10166 127410 10218
rect 127410 10166 127412 10218
rect 127356 10164 127412 10166
rect 127460 10218 127516 10220
rect 127460 10166 127462 10218
rect 127462 10166 127514 10218
rect 127514 10166 127516 10218
rect 127460 10164 127516 10166
rect 127564 10218 127620 10220
rect 127564 10166 127566 10218
rect 127566 10166 127618 10218
rect 127618 10166 127620 10218
rect 127564 10164 127620 10166
rect 158076 10218 158132 10220
rect 158076 10166 158078 10218
rect 158078 10166 158130 10218
rect 158130 10166 158132 10218
rect 158076 10164 158132 10166
rect 158180 10218 158236 10220
rect 158180 10166 158182 10218
rect 158182 10166 158234 10218
rect 158234 10166 158236 10218
rect 158180 10164 158236 10166
rect 158284 10218 158340 10220
rect 158284 10166 158286 10218
rect 158286 10166 158338 10218
rect 158338 10166 158340 10218
rect 158284 10164 158340 10166
rect 188796 10218 188852 10220
rect 188796 10166 188798 10218
rect 188798 10166 188850 10218
rect 188850 10166 188852 10218
rect 188796 10164 188852 10166
rect 188900 10218 188956 10220
rect 188900 10166 188902 10218
rect 188902 10166 188954 10218
rect 188954 10166 188956 10218
rect 188900 10164 188956 10166
rect 189004 10218 189060 10220
rect 189004 10166 189006 10218
rect 189006 10166 189058 10218
rect 189058 10166 189060 10218
rect 189004 10164 189060 10166
rect 12684 9548 12740 9604
rect 2492 9436 2548 9492
rect 5136 9434 5192 9436
rect 5136 9382 5138 9434
rect 5138 9382 5190 9434
rect 5190 9382 5192 9434
rect 5136 9380 5192 9382
rect 5240 9434 5296 9436
rect 5240 9382 5242 9434
rect 5242 9382 5294 9434
rect 5294 9382 5296 9434
rect 5240 9380 5296 9382
rect 5344 9434 5400 9436
rect 5344 9382 5346 9434
rect 5346 9382 5398 9434
rect 5398 9382 5400 9434
rect 5344 9380 5400 9382
rect 35856 9434 35912 9436
rect 35856 9382 35858 9434
rect 35858 9382 35910 9434
rect 35910 9382 35912 9434
rect 35856 9380 35912 9382
rect 35960 9434 36016 9436
rect 35960 9382 35962 9434
rect 35962 9382 36014 9434
rect 36014 9382 36016 9434
rect 35960 9380 36016 9382
rect 36064 9434 36120 9436
rect 36064 9382 36066 9434
rect 36066 9382 36118 9434
rect 36118 9382 36120 9434
rect 36064 9380 36120 9382
rect 66576 9434 66632 9436
rect 66576 9382 66578 9434
rect 66578 9382 66630 9434
rect 66630 9382 66632 9434
rect 66576 9380 66632 9382
rect 66680 9434 66736 9436
rect 66680 9382 66682 9434
rect 66682 9382 66734 9434
rect 66734 9382 66736 9434
rect 66680 9380 66736 9382
rect 66784 9434 66840 9436
rect 66784 9382 66786 9434
rect 66786 9382 66838 9434
rect 66838 9382 66840 9434
rect 66784 9380 66840 9382
rect 97296 9434 97352 9436
rect 97296 9382 97298 9434
rect 97298 9382 97350 9434
rect 97350 9382 97352 9434
rect 97296 9380 97352 9382
rect 97400 9434 97456 9436
rect 97400 9382 97402 9434
rect 97402 9382 97454 9434
rect 97454 9382 97456 9434
rect 97400 9380 97456 9382
rect 97504 9434 97560 9436
rect 97504 9382 97506 9434
rect 97506 9382 97558 9434
rect 97558 9382 97560 9434
rect 97504 9380 97560 9382
rect 128016 9434 128072 9436
rect 128016 9382 128018 9434
rect 128018 9382 128070 9434
rect 128070 9382 128072 9434
rect 128016 9380 128072 9382
rect 128120 9434 128176 9436
rect 128120 9382 128122 9434
rect 128122 9382 128174 9434
rect 128174 9382 128176 9434
rect 128120 9380 128176 9382
rect 128224 9434 128280 9436
rect 128224 9382 128226 9434
rect 128226 9382 128278 9434
rect 128278 9382 128280 9434
rect 128224 9380 128280 9382
rect 158736 9434 158792 9436
rect 158736 9382 158738 9434
rect 158738 9382 158790 9434
rect 158790 9382 158792 9434
rect 158736 9380 158792 9382
rect 158840 9434 158896 9436
rect 158840 9382 158842 9434
rect 158842 9382 158894 9434
rect 158894 9382 158896 9434
rect 158840 9380 158896 9382
rect 158944 9434 159000 9436
rect 158944 9382 158946 9434
rect 158946 9382 158998 9434
rect 158998 9382 159000 9434
rect 158944 9380 159000 9382
rect 189456 9434 189512 9436
rect 189456 9382 189458 9434
rect 189458 9382 189510 9434
rect 189510 9382 189512 9434
rect 189456 9380 189512 9382
rect 189560 9434 189616 9436
rect 189560 9382 189562 9434
rect 189562 9382 189614 9434
rect 189614 9382 189616 9434
rect 189560 9380 189616 9382
rect 189664 9434 189720 9436
rect 189664 9382 189666 9434
rect 189666 9382 189718 9434
rect 189718 9382 189720 9434
rect 189664 9380 189720 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 127356 8650 127412 8652
rect 127356 8598 127358 8650
rect 127358 8598 127410 8650
rect 127410 8598 127412 8650
rect 127356 8596 127412 8598
rect 127460 8650 127516 8652
rect 127460 8598 127462 8650
rect 127462 8598 127514 8650
rect 127514 8598 127516 8650
rect 127460 8596 127516 8598
rect 127564 8650 127620 8652
rect 127564 8598 127566 8650
rect 127566 8598 127618 8650
rect 127618 8598 127620 8650
rect 127564 8596 127620 8598
rect 158076 8650 158132 8652
rect 158076 8598 158078 8650
rect 158078 8598 158130 8650
rect 158130 8598 158132 8650
rect 158076 8596 158132 8598
rect 158180 8650 158236 8652
rect 158180 8598 158182 8650
rect 158182 8598 158234 8650
rect 158234 8598 158236 8650
rect 158180 8596 158236 8598
rect 158284 8650 158340 8652
rect 158284 8598 158286 8650
rect 158286 8598 158338 8650
rect 158338 8598 158340 8650
rect 158284 8596 158340 8598
rect 188796 8650 188852 8652
rect 188796 8598 188798 8650
rect 188798 8598 188850 8650
rect 188850 8598 188852 8650
rect 188796 8596 188852 8598
rect 188900 8650 188956 8652
rect 188900 8598 188902 8650
rect 188902 8598 188954 8650
rect 188954 8598 188956 8650
rect 188900 8596 188956 8598
rect 189004 8650 189060 8652
rect 189004 8598 189006 8650
rect 189006 8598 189058 8650
rect 189058 8598 189060 8650
rect 189004 8596 189060 8598
rect 5136 7866 5192 7868
rect 5136 7814 5138 7866
rect 5138 7814 5190 7866
rect 5190 7814 5192 7866
rect 5136 7812 5192 7814
rect 5240 7866 5296 7868
rect 5240 7814 5242 7866
rect 5242 7814 5294 7866
rect 5294 7814 5296 7866
rect 5240 7812 5296 7814
rect 5344 7866 5400 7868
rect 5344 7814 5346 7866
rect 5346 7814 5398 7866
rect 5398 7814 5400 7866
rect 5344 7812 5400 7814
rect 35856 7866 35912 7868
rect 35856 7814 35858 7866
rect 35858 7814 35910 7866
rect 35910 7814 35912 7866
rect 35856 7812 35912 7814
rect 35960 7866 36016 7868
rect 35960 7814 35962 7866
rect 35962 7814 36014 7866
rect 36014 7814 36016 7866
rect 35960 7812 36016 7814
rect 36064 7866 36120 7868
rect 36064 7814 36066 7866
rect 36066 7814 36118 7866
rect 36118 7814 36120 7866
rect 36064 7812 36120 7814
rect 66576 7866 66632 7868
rect 66576 7814 66578 7866
rect 66578 7814 66630 7866
rect 66630 7814 66632 7866
rect 66576 7812 66632 7814
rect 66680 7866 66736 7868
rect 66680 7814 66682 7866
rect 66682 7814 66734 7866
rect 66734 7814 66736 7866
rect 66680 7812 66736 7814
rect 66784 7866 66840 7868
rect 66784 7814 66786 7866
rect 66786 7814 66838 7866
rect 66838 7814 66840 7866
rect 66784 7812 66840 7814
rect 97296 7866 97352 7868
rect 97296 7814 97298 7866
rect 97298 7814 97350 7866
rect 97350 7814 97352 7866
rect 97296 7812 97352 7814
rect 97400 7866 97456 7868
rect 97400 7814 97402 7866
rect 97402 7814 97454 7866
rect 97454 7814 97456 7866
rect 97400 7812 97456 7814
rect 97504 7866 97560 7868
rect 97504 7814 97506 7866
rect 97506 7814 97558 7866
rect 97558 7814 97560 7866
rect 97504 7812 97560 7814
rect 128016 7866 128072 7868
rect 128016 7814 128018 7866
rect 128018 7814 128070 7866
rect 128070 7814 128072 7866
rect 128016 7812 128072 7814
rect 128120 7866 128176 7868
rect 128120 7814 128122 7866
rect 128122 7814 128174 7866
rect 128174 7814 128176 7866
rect 128120 7812 128176 7814
rect 128224 7866 128280 7868
rect 128224 7814 128226 7866
rect 128226 7814 128278 7866
rect 128278 7814 128280 7866
rect 128224 7812 128280 7814
rect 158736 7866 158792 7868
rect 158736 7814 158738 7866
rect 158738 7814 158790 7866
rect 158790 7814 158792 7866
rect 158736 7812 158792 7814
rect 158840 7866 158896 7868
rect 158840 7814 158842 7866
rect 158842 7814 158894 7866
rect 158894 7814 158896 7866
rect 158840 7812 158896 7814
rect 158944 7866 159000 7868
rect 158944 7814 158946 7866
rect 158946 7814 158998 7866
rect 158998 7814 159000 7866
rect 158944 7812 159000 7814
rect 189456 7866 189512 7868
rect 189456 7814 189458 7866
rect 189458 7814 189510 7866
rect 189510 7814 189512 7866
rect 189456 7812 189512 7814
rect 189560 7866 189616 7868
rect 189560 7814 189562 7866
rect 189562 7814 189614 7866
rect 189614 7814 189616 7866
rect 189560 7812 189616 7814
rect 189664 7866 189720 7868
rect 189664 7814 189666 7866
rect 189666 7814 189718 7866
rect 189718 7814 189720 7866
rect 189664 7812 189720 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 127356 7082 127412 7084
rect 127356 7030 127358 7082
rect 127358 7030 127410 7082
rect 127410 7030 127412 7082
rect 127356 7028 127412 7030
rect 127460 7082 127516 7084
rect 127460 7030 127462 7082
rect 127462 7030 127514 7082
rect 127514 7030 127516 7082
rect 127460 7028 127516 7030
rect 127564 7082 127620 7084
rect 127564 7030 127566 7082
rect 127566 7030 127618 7082
rect 127618 7030 127620 7082
rect 127564 7028 127620 7030
rect 158076 7082 158132 7084
rect 158076 7030 158078 7082
rect 158078 7030 158130 7082
rect 158130 7030 158132 7082
rect 158076 7028 158132 7030
rect 158180 7082 158236 7084
rect 158180 7030 158182 7082
rect 158182 7030 158234 7082
rect 158234 7030 158236 7082
rect 158180 7028 158236 7030
rect 158284 7082 158340 7084
rect 158284 7030 158286 7082
rect 158286 7030 158338 7082
rect 158338 7030 158340 7082
rect 158284 7028 158340 7030
rect 188796 7082 188852 7084
rect 188796 7030 188798 7082
rect 188798 7030 188850 7082
rect 188850 7030 188852 7082
rect 188796 7028 188852 7030
rect 188900 7082 188956 7084
rect 188900 7030 188902 7082
rect 188902 7030 188954 7082
rect 188954 7030 188956 7082
rect 188900 7028 188956 7030
rect 189004 7082 189060 7084
rect 189004 7030 189006 7082
rect 189006 7030 189058 7082
rect 189058 7030 189060 7082
rect 189004 7028 189060 7030
rect 5136 6298 5192 6300
rect 5136 6246 5138 6298
rect 5138 6246 5190 6298
rect 5190 6246 5192 6298
rect 5136 6244 5192 6246
rect 5240 6298 5296 6300
rect 5240 6246 5242 6298
rect 5242 6246 5294 6298
rect 5294 6246 5296 6298
rect 5240 6244 5296 6246
rect 5344 6298 5400 6300
rect 5344 6246 5346 6298
rect 5346 6246 5398 6298
rect 5398 6246 5400 6298
rect 5344 6244 5400 6246
rect 35856 6298 35912 6300
rect 35856 6246 35858 6298
rect 35858 6246 35910 6298
rect 35910 6246 35912 6298
rect 35856 6244 35912 6246
rect 35960 6298 36016 6300
rect 35960 6246 35962 6298
rect 35962 6246 36014 6298
rect 36014 6246 36016 6298
rect 35960 6244 36016 6246
rect 36064 6298 36120 6300
rect 36064 6246 36066 6298
rect 36066 6246 36118 6298
rect 36118 6246 36120 6298
rect 36064 6244 36120 6246
rect 66576 6298 66632 6300
rect 66576 6246 66578 6298
rect 66578 6246 66630 6298
rect 66630 6246 66632 6298
rect 66576 6244 66632 6246
rect 66680 6298 66736 6300
rect 66680 6246 66682 6298
rect 66682 6246 66734 6298
rect 66734 6246 66736 6298
rect 66680 6244 66736 6246
rect 66784 6298 66840 6300
rect 66784 6246 66786 6298
rect 66786 6246 66838 6298
rect 66838 6246 66840 6298
rect 66784 6244 66840 6246
rect 97296 6298 97352 6300
rect 97296 6246 97298 6298
rect 97298 6246 97350 6298
rect 97350 6246 97352 6298
rect 97296 6244 97352 6246
rect 97400 6298 97456 6300
rect 97400 6246 97402 6298
rect 97402 6246 97454 6298
rect 97454 6246 97456 6298
rect 97400 6244 97456 6246
rect 97504 6298 97560 6300
rect 97504 6246 97506 6298
rect 97506 6246 97558 6298
rect 97558 6246 97560 6298
rect 97504 6244 97560 6246
rect 128016 6298 128072 6300
rect 128016 6246 128018 6298
rect 128018 6246 128070 6298
rect 128070 6246 128072 6298
rect 128016 6244 128072 6246
rect 128120 6298 128176 6300
rect 128120 6246 128122 6298
rect 128122 6246 128174 6298
rect 128174 6246 128176 6298
rect 128120 6244 128176 6246
rect 128224 6298 128280 6300
rect 128224 6246 128226 6298
rect 128226 6246 128278 6298
rect 128278 6246 128280 6298
rect 128224 6244 128280 6246
rect 158736 6298 158792 6300
rect 158736 6246 158738 6298
rect 158738 6246 158790 6298
rect 158790 6246 158792 6298
rect 158736 6244 158792 6246
rect 158840 6298 158896 6300
rect 158840 6246 158842 6298
rect 158842 6246 158894 6298
rect 158894 6246 158896 6298
rect 158840 6244 158896 6246
rect 158944 6298 159000 6300
rect 158944 6246 158946 6298
rect 158946 6246 158998 6298
rect 158998 6246 159000 6298
rect 158944 6244 159000 6246
rect 189456 6298 189512 6300
rect 189456 6246 189458 6298
rect 189458 6246 189510 6298
rect 189510 6246 189512 6298
rect 189456 6244 189512 6246
rect 189560 6298 189616 6300
rect 189560 6246 189562 6298
rect 189562 6246 189614 6298
rect 189614 6246 189616 6298
rect 189560 6244 189616 6246
rect 189664 6298 189720 6300
rect 189664 6246 189666 6298
rect 189666 6246 189718 6298
rect 189718 6246 189720 6298
rect 189664 6244 189720 6246
rect 1708 5628 1764 5684
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 127356 5514 127412 5516
rect 127356 5462 127358 5514
rect 127358 5462 127410 5514
rect 127410 5462 127412 5514
rect 127356 5460 127412 5462
rect 127460 5514 127516 5516
rect 127460 5462 127462 5514
rect 127462 5462 127514 5514
rect 127514 5462 127516 5514
rect 127460 5460 127516 5462
rect 127564 5514 127620 5516
rect 127564 5462 127566 5514
rect 127566 5462 127618 5514
rect 127618 5462 127620 5514
rect 127564 5460 127620 5462
rect 158076 5514 158132 5516
rect 158076 5462 158078 5514
rect 158078 5462 158130 5514
rect 158130 5462 158132 5514
rect 158076 5460 158132 5462
rect 158180 5514 158236 5516
rect 158180 5462 158182 5514
rect 158182 5462 158234 5514
rect 158234 5462 158236 5514
rect 158180 5460 158236 5462
rect 158284 5514 158340 5516
rect 158284 5462 158286 5514
rect 158286 5462 158338 5514
rect 158338 5462 158340 5514
rect 158284 5460 158340 5462
rect 188796 5514 188852 5516
rect 188796 5462 188798 5514
rect 188798 5462 188850 5514
rect 188850 5462 188852 5514
rect 188796 5460 188852 5462
rect 188900 5514 188956 5516
rect 188900 5462 188902 5514
rect 188902 5462 188954 5514
rect 188954 5462 188956 5514
rect 188900 5460 188956 5462
rect 189004 5514 189060 5516
rect 189004 5462 189006 5514
rect 189006 5462 189058 5514
rect 189058 5462 189060 5514
rect 189004 5460 189060 5462
rect 5136 4730 5192 4732
rect 5136 4678 5138 4730
rect 5138 4678 5190 4730
rect 5190 4678 5192 4730
rect 5136 4676 5192 4678
rect 5240 4730 5296 4732
rect 5240 4678 5242 4730
rect 5242 4678 5294 4730
rect 5294 4678 5296 4730
rect 5240 4676 5296 4678
rect 5344 4730 5400 4732
rect 5344 4678 5346 4730
rect 5346 4678 5398 4730
rect 5398 4678 5400 4730
rect 5344 4676 5400 4678
rect 35856 4730 35912 4732
rect 35856 4678 35858 4730
rect 35858 4678 35910 4730
rect 35910 4678 35912 4730
rect 35856 4676 35912 4678
rect 35960 4730 36016 4732
rect 35960 4678 35962 4730
rect 35962 4678 36014 4730
rect 36014 4678 36016 4730
rect 35960 4676 36016 4678
rect 36064 4730 36120 4732
rect 36064 4678 36066 4730
rect 36066 4678 36118 4730
rect 36118 4678 36120 4730
rect 36064 4676 36120 4678
rect 66576 4730 66632 4732
rect 66576 4678 66578 4730
rect 66578 4678 66630 4730
rect 66630 4678 66632 4730
rect 66576 4676 66632 4678
rect 66680 4730 66736 4732
rect 66680 4678 66682 4730
rect 66682 4678 66734 4730
rect 66734 4678 66736 4730
rect 66680 4676 66736 4678
rect 66784 4730 66840 4732
rect 66784 4678 66786 4730
rect 66786 4678 66838 4730
rect 66838 4678 66840 4730
rect 66784 4676 66840 4678
rect 97296 4730 97352 4732
rect 97296 4678 97298 4730
rect 97298 4678 97350 4730
rect 97350 4678 97352 4730
rect 97296 4676 97352 4678
rect 97400 4730 97456 4732
rect 97400 4678 97402 4730
rect 97402 4678 97454 4730
rect 97454 4678 97456 4730
rect 97400 4676 97456 4678
rect 97504 4730 97560 4732
rect 97504 4678 97506 4730
rect 97506 4678 97558 4730
rect 97558 4678 97560 4730
rect 97504 4676 97560 4678
rect 128016 4730 128072 4732
rect 128016 4678 128018 4730
rect 128018 4678 128070 4730
rect 128070 4678 128072 4730
rect 128016 4676 128072 4678
rect 128120 4730 128176 4732
rect 128120 4678 128122 4730
rect 128122 4678 128174 4730
rect 128174 4678 128176 4730
rect 128120 4676 128176 4678
rect 128224 4730 128280 4732
rect 128224 4678 128226 4730
rect 128226 4678 128278 4730
rect 128278 4678 128280 4730
rect 128224 4676 128280 4678
rect 158736 4730 158792 4732
rect 158736 4678 158738 4730
rect 158738 4678 158790 4730
rect 158790 4678 158792 4730
rect 158736 4676 158792 4678
rect 158840 4730 158896 4732
rect 158840 4678 158842 4730
rect 158842 4678 158894 4730
rect 158894 4678 158896 4730
rect 158840 4676 158896 4678
rect 158944 4730 159000 4732
rect 158944 4678 158946 4730
rect 158946 4678 158998 4730
rect 158998 4678 159000 4730
rect 158944 4676 159000 4678
rect 189456 4730 189512 4732
rect 189456 4678 189458 4730
rect 189458 4678 189510 4730
rect 189510 4678 189512 4730
rect 189456 4676 189512 4678
rect 189560 4730 189616 4732
rect 189560 4678 189562 4730
rect 189562 4678 189614 4730
rect 189614 4678 189616 4730
rect 189560 4676 189616 4678
rect 189664 4730 189720 4732
rect 189664 4678 189666 4730
rect 189666 4678 189718 4730
rect 189718 4678 189720 4730
rect 189664 4676 189720 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 127356 3946 127412 3948
rect 127356 3894 127358 3946
rect 127358 3894 127410 3946
rect 127410 3894 127412 3946
rect 127356 3892 127412 3894
rect 127460 3946 127516 3948
rect 127460 3894 127462 3946
rect 127462 3894 127514 3946
rect 127514 3894 127516 3946
rect 127460 3892 127516 3894
rect 127564 3946 127620 3948
rect 127564 3894 127566 3946
rect 127566 3894 127618 3946
rect 127618 3894 127620 3946
rect 127564 3892 127620 3894
rect 158076 3946 158132 3948
rect 158076 3894 158078 3946
rect 158078 3894 158130 3946
rect 158130 3894 158132 3946
rect 158076 3892 158132 3894
rect 158180 3946 158236 3948
rect 158180 3894 158182 3946
rect 158182 3894 158234 3946
rect 158234 3894 158236 3946
rect 158180 3892 158236 3894
rect 158284 3946 158340 3948
rect 158284 3894 158286 3946
rect 158286 3894 158338 3946
rect 158338 3894 158340 3946
rect 158284 3892 158340 3894
rect 188796 3946 188852 3948
rect 188796 3894 188798 3946
rect 188798 3894 188850 3946
rect 188850 3894 188852 3946
rect 188796 3892 188852 3894
rect 188900 3946 188956 3948
rect 188900 3894 188902 3946
rect 188902 3894 188954 3946
rect 188954 3894 188956 3946
rect 188900 3892 188956 3894
rect 189004 3946 189060 3948
rect 189004 3894 189006 3946
rect 189006 3894 189058 3946
rect 189058 3894 189060 3946
rect 189004 3892 189060 3894
rect 5136 3162 5192 3164
rect 5136 3110 5138 3162
rect 5138 3110 5190 3162
rect 5190 3110 5192 3162
rect 5136 3108 5192 3110
rect 5240 3162 5296 3164
rect 5240 3110 5242 3162
rect 5242 3110 5294 3162
rect 5294 3110 5296 3162
rect 5240 3108 5296 3110
rect 5344 3162 5400 3164
rect 5344 3110 5346 3162
rect 5346 3110 5398 3162
rect 5398 3110 5400 3162
rect 5344 3108 5400 3110
rect 1708 1820 1764 1876
rect 35856 3162 35912 3164
rect 35856 3110 35858 3162
rect 35858 3110 35910 3162
rect 35910 3110 35912 3162
rect 35856 3108 35912 3110
rect 35960 3162 36016 3164
rect 35960 3110 35962 3162
rect 35962 3110 36014 3162
rect 36014 3110 36016 3162
rect 35960 3108 36016 3110
rect 36064 3162 36120 3164
rect 36064 3110 36066 3162
rect 36066 3110 36118 3162
rect 36118 3110 36120 3162
rect 36064 3108 36120 3110
rect 66576 3162 66632 3164
rect 66576 3110 66578 3162
rect 66578 3110 66630 3162
rect 66630 3110 66632 3162
rect 66576 3108 66632 3110
rect 66680 3162 66736 3164
rect 66680 3110 66682 3162
rect 66682 3110 66734 3162
rect 66734 3110 66736 3162
rect 66680 3108 66736 3110
rect 66784 3162 66840 3164
rect 66784 3110 66786 3162
rect 66786 3110 66838 3162
rect 66838 3110 66840 3162
rect 66784 3108 66840 3110
rect 97296 3162 97352 3164
rect 97296 3110 97298 3162
rect 97298 3110 97350 3162
rect 97350 3110 97352 3162
rect 97296 3108 97352 3110
rect 97400 3162 97456 3164
rect 97400 3110 97402 3162
rect 97402 3110 97454 3162
rect 97454 3110 97456 3162
rect 97400 3108 97456 3110
rect 97504 3162 97560 3164
rect 97504 3110 97506 3162
rect 97506 3110 97558 3162
rect 97558 3110 97560 3162
rect 97504 3108 97560 3110
rect 128016 3162 128072 3164
rect 128016 3110 128018 3162
rect 128018 3110 128070 3162
rect 128070 3110 128072 3162
rect 128016 3108 128072 3110
rect 128120 3162 128176 3164
rect 128120 3110 128122 3162
rect 128122 3110 128174 3162
rect 128174 3110 128176 3162
rect 128120 3108 128176 3110
rect 128224 3162 128280 3164
rect 128224 3110 128226 3162
rect 128226 3110 128278 3162
rect 128278 3110 128280 3162
rect 128224 3108 128280 3110
rect 158736 3162 158792 3164
rect 158736 3110 158738 3162
rect 158738 3110 158790 3162
rect 158790 3110 158792 3162
rect 158736 3108 158792 3110
rect 158840 3162 158896 3164
rect 158840 3110 158842 3162
rect 158842 3110 158894 3162
rect 158894 3110 158896 3162
rect 158840 3108 158896 3110
rect 158944 3162 159000 3164
rect 158944 3110 158946 3162
rect 158946 3110 158998 3162
rect 158998 3110 159000 3162
rect 158944 3108 159000 3110
rect 189456 3162 189512 3164
rect 189456 3110 189458 3162
rect 189458 3110 189510 3162
rect 189510 3110 189512 3162
rect 189456 3108 189512 3110
rect 189560 3162 189616 3164
rect 189560 3110 189562 3162
rect 189562 3110 189614 3162
rect 189614 3110 189616 3162
rect 189560 3108 189616 3110
rect 189664 3162 189720 3164
rect 189664 3110 189666 3162
rect 189666 3110 189718 3162
rect 189718 3110 189720 3162
rect 189664 3108 189720 3110
<< metal3 >>
rect 0 158004 800 158032
rect 0 157948 1764 158004
rect 0 157920 800 157948
rect 1708 157892 1764 157948
rect 1698 157836 1708 157892
rect 1764 157836 1774 157892
rect 5126 156772 5136 156828
rect 5192 156772 5240 156828
rect 5296 156772 5344 156828
rect 5400 156772 5410 156828
rect 35846 156772 35856 156828
rect 35912 156772 35960 156828
rect 36016 156772 36064 156828
rect 36120 156772 36130 156828
rect 66566 156772 66576 156828
rect 66632 156772 66680 156828
rect 66736 156772 66784 156828
rect 66840 156772 66850 156828
rect 97286 156772 97296 156828
rect 97352 156772 97400 156828
rect 97456 156772 97504 156828
rect 97560 156772 97570 156828
rect 128006 156772 128016 156828
rect 128072 156772 128120 156828
rect 128176 156772 128224 156828
rect 128280 156772 128290 156828
rect 158726 156772 158736 156828
rect 158792 156772 158840 156828
rect 158896 156772 158944 156828
rect 159000 156772 159010 156828
rect 189446 156772 189456 156828
rect 189512 156772 189560 156828
rect 189616 156772 189664 156828
rect 189720 156772 189730 156828
rect 41906 156604 41916 156660
rect 41972 156604 43708 156660
rect 43764 156604 43774 156660
rect 64754 156604 64764 156660
rect 64820 156604 66556 156660
rect 66612 156604 66622 156660
rect 134194 156604 134204 156660
rect 134260 156604 135100 156660
rect 135156 156604 135166 156660
rect 63746 156492 63756 156548
rect 63812 156492 87612 156548
rect 87668 156492 87678 156548
rect 65090 156380 65100 156436
rect 65156 156380 67228 156436
rect 67172 156324 67228 156380
rect 20066 156268 20076 156324
rect 20132 156268 22764 156324
rect 22820 156268 22830 156324
rect 42802 156268 42812 156324
rect 42868 156268 56252 156324
rect 56308 156268 56318 156324
rect 64418 156268 64428 156324
rect 64484 156268 65324 156324
rect 65380 156268 65390 156324
rect 67172 156268 111132 156324
rect 111188 156268 111198 156324
rect 4466 155988 4476 156044
rect 4532 155988 4580 156044
rect 4636 155988 4684 156044
rect 4740 155988 4750 156044
rect 35186 155988 35196 156044
rect 35252 155988 35300 156044
rect 35356 155988 35404 156044
rect 35460 155988 35470 156044
rect 65906 155988 65916 156044
rect 65972 155988 66020 156044
rect 66076 155988 66124 156044
rect 66180 155988 66190 156044
rect 96626 155988 96636 156044
rect 96692 155988 96740 156044
rect 96796 155988 96844 156044
rect 96900 155988 96910 156044
rect 127346 155988 127356 156044
rect 127412 155988 127460 156044
rect 127516 155988 127564 156044
rect 127620 155988 127630 156044
rect 158066 155988 158076 156044
rect 158132 155988 158180 156044
rect 158236 155988 158284 156044
rect 158340 155988 158350 156044
rect 188786 155988 188796 156044
rect 188852 155988 188900 156044
rect 188956 155988 189004 156044
rect 189060 155988 189070 156044
rect 194226 155820 194236 155876
rect 194292 155820 194908 155876
rect 194964 155820 194974 155876
rect 5126 155204 5136 155260
rect 5192 155204 5240 155260
rect 5296 155204 5344 155260
rect 5400 155204 5410 155260
rect 35846 155204 35856 155260
rect 35912 155204 35960 155260
rect 36016 155204 36064 155260
rect 36120 155204 36130 155260
rect 66566 155204 66576 155260
rect 66632 155204 66680 155260
rect 66736 155204 66784 155260
rect 66840 155204 66850 155260
rect 97286 155204 97296 155260
rect 97352 155204 97400 155260
rect 97456 155204 97504 155260
rect 97560 155204 97570 155260
rect 128006 155204 128016 155260
rect 128072 155204 128120 155260
rect 128176 155204 128224 155260
rect 128280 155204 128290 155260
rect 158726 155204 158736 155260
rect 158792 155204 158840 155260
rect 158896 155204 158944 155260
rect 159000 155204 159010 155260
rect 189446 155204 189456 155260
rect 189512 155204 189560 155260
rect 189616 155204 189664 155260
rect 189720 155204 189730 155260
rect 4466 154420 4476 154476
rect 4532 154420 4580 154476
rect 4636 154420 4684 154476
rect 4740 154420 4750 154476
rect 35186 154420 35196 154476
rect 35252 154420 35300 154476
rect 35356 154420 35404 154476
rect 35460 154420 35470 154476
rect 65906 154420 65916 154476
rect 65972 154420 66020 154476
rect 66076 154420 66124 154476
rect 66180 154420 66190 154476
rect 96626 154420 96636 154476
rect 96692 154420 96740 154476
rect 96796 154420 96844 154476
rect 96900 154420 96910 154476
rect 127346 154420 127356 154476
rect 127412 154420 127460 154476
rect 127516 154420 127564 154476
rect 127620 154420 127630 154476
rect 158066 154420 158076 154476
rect 158132 154420 158180 154476
rect 158236 154420 158284 154476
rect 158340 154420 158350 154476
rect 188786 154420 188796 154476
rect 188852 154420 188900 154476
rect 188956 154420 189004 154476
rect 189060 154420 189070 154476
rect 0 154196 800 154224
rect 205332 154196 206132 154224
rect 0 154140 1708 154196
rect 1764 154140 1774 154196
rect 204306 154140 204316 154196
rect 204372 154140 206132 154196
rect 0 154112 800 154140
rect 205332 154112 206132 154140
rect 5126 153636 5136 153692
rect 5192 153636 5240 153692
rect 5296 153636 5344 153692
rect 5400 153636 5410 153692
rect 35846 153636 35856 153692
rect 35912 153636 35960 153692
rect 36016 153636 36064 153692
rect 36120 153636 36130 153692
rect 66566 153636 66576 153692
rect 66632 153636 66680 153692
rect 66736 153636 66784 153692
rect 66840 153636 66850 153692
rect 97286 153636 97296 153692
rect 97352 153636 97400 153692
rect 97456 153636 97504 153692
rect 97560 153636 97570 153692
rect 128006 153636 128016 153692
rect 128072 153636 128120 153692
rect 128176 153636 128224 153692
rect 128280 153636 128290 153692
rect 158726 153636 158736 153692
rect 158792 153636 158840 153692
rect 158896 153636 158944 153692
rect 159000 153636 159010 153692
rect 189446 153636 189456 153692
rect 189512 153636 189560 153692
rect 189616 153636 189664 153692
rect 189720 153636 189730 153692
rect 4466 152852 4476 152908
rect 4532 152852 4580 152908
rect 4636 152852 4684 152908
rect 4740 152852 4750 152908
rect 35186 152852 35196 152908
rect 35252 152852 35300 152908
rect 35356 152852 35404 152908
rect 35460 152852 35470 152908
rect 65906 152852 65916 152908
rect 65972 152852 66020 152908
rect 66076 152852 66124 152908
rect 66180 152852 66190 152908
rect 96626 152852 96636 152908
rect 96692 152852 96740 152908
rect 96796 152852 96844 152908
rect 96900 152852 96910 152908
rect 127346 152852 127356 152908
rect 127412 152852 127460 152908
rect 127516 152852 127564 152908
rect 127620 152852 127630 152908
rect 158066 152852 158076 152908
rect 158132 152852 158180 152908
rect 158236 152852 158284 152908
rect 158340 152852 158350 152908
rect 188786 152852 188796 152908
rect 188852 152852 188900 152908
rect 188956 152852 189004 152908
rect 189060 152852 189070 152908
rect 5126 152068 5136 152124
rect 5192 152068 5240 152124
rect 5296 152068 5344 152124
rect 5400 152068 5410 152124
rect 35846 152068 35856 152124
rect 35912 152068 35960 152124
rect 36016 152068 36064 152124
rect 36120 152068 36130 152124
rect 66566 152068 66576 152124
rect 66632 152068 66680 152124
rect 66736 152068 66784 152124
rect 66840 152068 66850 152124
rect 97286 152068 97296 152124
rect 97352 152068 97400 152124
rect 97456 152068 97504 152124
rect 97560 152068 97570 152124
rect 128006 152068 128016 152124
rect 128072 152068 128120 152124
rect 128176 152068 128224 152124
rect 128280 152068 128290 152124
rect 158726 152068 158736 152124
rect 158792 152068 158840 152124
rect 158896 152068 158944 152124
rect 159000 152068 159010 152124
rect 189446 152068 189456 152124
rect 189512 152068 189560 152124
rect 189616 152068 189664 152124
rect 189720 152068 189730 152124
rect 4466 151284 4476 151340
rect 4532 151284 4580 151340
rect 4636 151284 4684 151340
rect 4740 151284 4750 151340
rect 35186 151284 35196 151340
rect 35252 151284 35300 151340
rect 35356 151284 35404 151340
rect 35460 151284 35470 151340
rect 65906 151284 65916 151340
rect 65972 151284 66020 151340
rect 66076 151284 66124 151340
rect 66180 151284 66190 151340
rect 96626 151284 96636 151340
rect 96692 151284 96740 151340
rect 96796 151284 96844 151340
rect 96900 151284 96910 151340
rect 127346 151284 127356 151340
rect 127412 151284 127460 151340
rect 127516 151284 127564 151340
rect 127620 151284 127630 151340
rect 158066 151284 158076 151340
rect 158132 151284 158180 151340
rect 158236 151284 158284 151340
rect 158340 151284 158350 151340
rect 188786 151284 188796 151340
rect 188852 151284 188900 151340
rect 188956 151284 189004 151340
rect 189060 151284 189070 151340
rect 5126 150500 5136 150556
rect 5192 150500 5240 150556
rect 5296 150500 5344 150556
rect 5400 150500 5410 150556
rect 35846 150500 35856 150556
rect 35912 150500 35960 150556
rect 36016 150500 36064 150556
rect 36120 150500 36130 150556
rect 66566 150500 66576 150556
rect 66632 150500 66680 150556
rect 66736 150500 66784 150556
rect 66840 150500 66850 150556
rect 97286 150500 97296 150556
rect 97352 150500 97400 150556
rect 97456 150500 97504 150556
rect 97560 150500 97570 150556
rect 128006 150500 128016 150556
rect 128072 150500 128120 150556
rect 128176 150500 128224 150556
rect 128280 150500 128290 150556
rect 158726 150500 158736 150556
rect 158792 150500 158840 150556
rect 158896 150500 158944 150556
rect 159000 150500 159010 150556
rect 189446 150500 189456 150556
rect 189512 150500 189560 150556
rect 189616 150500 189664 150556
rect 189720 150500 189730 150556
rect 0 150388 800 150416
rect 0 150332 1708 150388
rect 1764 150332 1774 150388
rect 0 150304 800 150332
rect 4466 149716 4476 149772
rect 4532 149716 4580 149772
rect 4636 149716 4684 149772
rect 4740 149716 4750 149772
rect 35186 149716 35196 149772
rect 35252 149716 35300 149772
rect 35356 149716 35404 149772
rect 35460 149716 35470 149772
rect 65906 149716 65916 149772
rect 65972 149716 66020 149772
rect 66076 149716 66124 149772
rect 66180 149716 66190 149772
rect 96626 149716 96636 149772
rect 96692 149716 96740 149772
rect 96796 149716 96844 149772
rect 96900 149716 96910 149772
rect 127346 149716 127356 149772
rect 127412 149716 127460 149772
rect 127516 149716 127564 149772
rect 127620 149716 127630 149772
rect 158066 149716 158076 149772
rect 158132 149716 158180 149772
rect 158236 149716 158284 149772
rect 158340 149716 158350 149772
rect 188786 149716 188796 149772
rect 188852 149716 188900 149772
rect 188956 149716 189004 149772
rect 189060 149716 189070 149772
rect 5126 148932 5136 148988
rect 5192 148932 5240 148988
rect 5296 148932 5344 148988
rect 5400 148932 5410 148988
rect 35846 148932 35856 148988
rect 35912 148932 35960 148988
rect 36016 148932 36064 148988
rect 36120 148932 36130 148988
rect 66566 148932 66576 148988
rect 66632 148932 66680 148988
rect 66736 148932 66784 148988
rect 66840 148932 66850 148988
rect 97286 148932 97296 148988
rect 97352 148932 97400 148988
rect 97456 148932 97504 148988
rect 97560 148932 97570 148988
rect 128006 148932 128016 148988
rect 128072 148932 128120 148988
rect 128176 148932 128224 148988
rect 128280 148932 128290 148988
rect 158726 148932 158736 148988
rect 158792 148932 158840 148988
rect 158896 148932 158944 148988
rect 159000 148932 159010 148988
rect 189446 148932 189456 148988
rect 189512 148932 189560 148988
rect 189616 148932 189664 148988
rect 189720 148932 189730 148988
rect 4466 148148 4476 148204
rect 4532 148148 4580 148204
rect 4636 148148 4684 148204
rect 4740 148148 4750 148204
rect 35186 148148 35196 148204
rect 35252 148148 35300 148204
rect 35356 148148 35404 148204
rect 35460 148148 35470 148204
rect 65906 148148 65916 148204
rect 65972 148148 66020 148204
rect 66076 148148 66124 148204
rect 66180 148148 66190 148204
rect 96626 148148 96636 148204
rect 96692 148148 96740 148204
rect 96796 148148 96844 148204
rect 96900 148148 96910 148204
rect 127346 148148 127356 148204
rect 127412 148148 127460 148204
rect 127516 148148 127564 148204
rect 127620 148148 127630 148204
rect 158066 148148 158076 148204
rect 158132 148148 158180 148204
rect 158236 148148 158284 148204
rect 158340 148148 158350 148204
rect 188786 148148 188796 148204
rect 188852 148148 188900 148204
rect 188956 148148 189004 148204
rect 189060 148148 189070 148204
rect 5126 147364 5136 147420
rect 5192 147364 5240 147420
rect 5296 147364 5344 147420
rect 5400 147364 5410 147420
rect 35846 147364 35856 147420
rect 35912 147364 35960 147420
rect 36016 147364 36064 147420
rect 36120 147364 36130 147420
rect 66566 147364 66576 147420
rect 66632 147364 66680 147420
rect 66736 147364 66784 147420
rect 66840 147364 66850 147420
rect 97286 147364 97296 147420
rect 97352 147364 97400 147420
rect 97456 147364 97504 147420
rect 97560 147364 97570 147420
rect 128006 147364 128016 147420
rect 128072 147364 128120 147420
rect 128176 147364 128224 147420
rect 128280 147364 128290 147420
rect 158726 147364 158736 147420
rect 158792 147364 158840 147420
rect 158896 147364 158944 147420
rect 159000 147364 159010 147420
rect 189446 147364 189456 147420
rect 189512 147364 189560 147420
rect 189616 147364 189664 147420
rect 189720 147364 189730 147420
rect 2818 146860 2828 146916
rect 2884 146860 12572 146916
rect 12628 146860 12638 146916
rect 0 146580 800 146608
rect 4466 146580 4476 146636
rect 4532 146580 4580 146636
rect 4636 146580 4684 146636
rect 4740 146580 4750 146636
rect 35186 146580 35196 146636
rect 35252 146580 35300 146636
rect 35356 146580 35404 146636
rect 35460 146580 35470 146636
rect 65906 146580 65916 146636
rect 65972 146580 66020 146636
rect 66076 146580 66124 146636
rect 66180 146580 66190 146636
rect 96626 146580 96636 146636
rect 96692 146580 96740 146636
rect 96796 146580 96844 146636
rect 96900 146580 96910 146636
rect 127346 146580 127356 146636
rect 127412 146580 127460 146636
rect 127516 146580 127564 146636
rect 127620 146580 127630 146636
rect 158066 146580 158076 146636
rect 158132 146580 158180 146636
rect 158236 146580 158284 146636
rect 158340 146580 158350 146636
rect 188786 146580 188796 146636
rect 188852 146580 188900 146636
rect 188956 146580 189004 146636
rect 189060 146580 189070 146636
rect 0 146524 1820 146580
rect 1876 146524 1886 146580
rect 0 146496 800 146524
rect 201058 146188 201068 146244
rect 201124 146188 201740 146244
rect 201796 146188 201806 146244
rect 5126 145796 5136 145852
rect 5192 145796 5240 145852
rect 5296 145796 5344 145852
rect 5400 145796 5410 145852
rect 35846 145796 35856 145852
rect 35912 145796 35960 145852
rect 36016 145796 36064 145852
rect 36120 145796 36130 145852
rect 66566 145796 66576 145852
rect 66632 145796 66680 145852
rect 66736 145796 66784 145852
rect 66840 145796 66850 145852
rect 97286 145796 97296 145852
rect 97352 145796 97400 145852
rect 97456 145796 97504 145852
rect 97560 145796 97570 145852
rect 128006 145796 128016 145852
rect 128072 145796 128120 145852
rect 128176 145796 128224 145852
rect 128280 145796 128290 145852
rect 158726 145796 158736 145852
rect 158792 145796 158840 145852
rect 158896 145796 158944 145852
rect 159000 145796 159010 145852
rect 189446 145796 189456 145852
rect 189512 145796 189560 145852
rect 189616 145796 189664 145852
rect 189720 145796 189730 145852
rect 205332 145460 206132 145488
rect 204082 145404 204092 145460
rect 204148 145404 206132 145460
rect 205332 145376 206132 145404
rect 4466 145012 4476 145068
rect 4532 145012 4580 145068
rect 4636 145012 4684 145068
rect 4740 145012 4750 145068
rect 35186 145012 35196 145068
rect 35252 145012 35300 145068
rect 35356 145012 35404 145068
rect 35460 145012 35470 145068
rect 65906 145012 65916 145068
rect 65972 145012 66020 145068
rect 66076 145012 66124 145068
rect 66180 145012 66190 145068
rect 96626 145012 96636 145068
rect 96692 145012 96740 145068
rect 96796 145012 96844 145068
rect 96900 145012 96910 145068
rect 127346 145012 127356 145068
rect 127412 145012 127460 145068
rect 127516 145012 127564 145068
rect 127620 145012 127630 145068
rect 158066 145012 158076 145068
rect 158132 145012 158180 145068
rect 158236 145012 158284 145068
rect 158340 145012 158350 145068
rect 188786 145012 188796 145068
rect 188852 145012 188900 145068
rect 188956 145012 189004 145068
rect 189060 145012 189070 145068
rect 5126 144228 5136 144284
rect 5192 144228 5240 144284
rect 5296 144228 5344 144284
rect 5400 144228 5410 144284
rect 189446 144228 189456 144284
rect 189512 144228 189560 144284
rect 189616 144228 189664 144284
rect 189720 144228 189730 144284
rect 4466 143444 4476 143500
rect 4532 143444 4580 143500
rect 4636 143444 4684 143500
rect 4740 143444 4750 143500
rect 188786 143444 188796 143500
rect 188852 143444 188900 143500
rect 188956 143444 189004 143500
rect 189060 143444 189070 143500
rect 0 142772 800 142800
rect 0 142716 1708 142772
rect 1764 142716 1774 142772
rect 0 142688 800 142716
rect 5126 142660 5136 142716
rect 5192 142660 5240 142716
rect 5296 142660 5344 142716
rect 5400 142660 5410 142716
rect 189446 142660 189456 142716
rect 189512 142660 189560 142716
rect 189616 142660 189664 142716
rect 189720 142660 189730 142716
rect 4466 141876 4476 141932
rect 4532 141876 4580 141932
rect 4636 141876 4684 141932
rect 4740 141876 4750 141932
rect 188786 141876 188796 141932
rect 188852 141876 188900 141932
rect 188956 141876 189004 141932
rect 189060 141876 189070 141932
rect 5126 141092 5136 141148
rect 5192 141092 5240 141148
rect 5296 141092 5344 141148
rect 5400 141092 5410 141148
rect 189446 141092 189456 141148
rect 189512 141092 189560 141148
rect 189616 141092 189664 141148
rect 189720 141092 189730 141148
rect 4466 140308 4476 140364
rect 4532 140308 4580 140364
rect 4636 140308 4684 140364
rect 4740 140308 4750 140364
rect 188786 140308 188796 140364
rect 188852 140308 188900 140364
rect 188956 140308 189004 140364
rect 189060 140308 189070 140364
rect 5126 139524 5136 139580
rect 5192 139524 5240 139580
rect 5296 139524 5344 139580
rect 5400 139524 5410 139580
rect 189446 139524 189456 139580
rect 189512 139524 189560 139580
rect 189616 139524 189664 139580
rect 189720 139524 189730 139580
rect 0 138964 800 138992
rect 0 138908 1708 138964
rect 1764 138908 1774 138964
rect 0 138880 800 138908
rect 4466 138740 4476 138796
rect 4532 138740 4580 138796
rect 4636 138740 4684 138796
rect 4740 138740 4750 138796
rect 188786 138740 188796 138796
rect 188852 138740 188900 138796
rect 188956 138740 189004 138796
rect 189060 138740 189070 138796
rect 5126 137956 5136 138012
rect 5192 137956 5240 138012
rect 5296 137956 5344 138012
rect 5400 137956 5410 138012
rect 189446 137956 189456 138012
rect 189512 137956 189560 138012
rect 189616 137956 189664 138012
rect 189720 137956 189730 138012
rect 4466 137172 4476 137228
rect 4532 137172 4580 137228
rect 4636 137172 4684 137228
rect 4740 137172 4750 137228
rect 188786 137172 188796 137228
rect 188852 137172 188900 137228
rect 188956 137172 189004 137228
rect 189060 137172 189070 137228
rect 205332 136640 206132 136752
rect 5126 136388 5136 136444
rect 5192 136388 5240 136444
rect 5296 136388 5344 136444
rect 5400 136388 5410 136444
rect 189446 136388 189456 136444
rect 189512 136388 189560 136444
rect 189616 136388 189664 136444
rect 189720 136388 189730 136444
rect 4466 135604 4476 135660
rect 4532 135604 4580 135660
rect 4636 135604 4684 135660
rect 4740 135604 4750 135660
rect 188786 135604 188796 135660
rect 188852 135604 188900 135660
rect 188956 135604 189004 135660
rect 189060 135604 189070 135660
rect 0 135156 800 135184
rect 0 135100 1708 135156
rect 1764 135100 1774 135156
rect 2818 135100 2828 135156
rect 2884 135100 17724 135156
rect 17780 135100 17790 135156
rect 0 135072 800 135100
rect 5126 134820 5136 134876
rect 5192 134820 5240 134876
rect 5296 134820 5344 134876
rect 5400 134820 5410 134876
rect 189446 134820 189456 134876
rect 189512 134820 189560 134876
rect 189616 134820 189664 134876
rect 189720 134820 189730 134876
rect 4466 134036 4476 134092
rect 4532 134036 4580 134092
rect 4636 134036 4684 134092
rect 4740 134036 4750 134092
rect 188786 134036 188796 134092
rect 188852 134036 188900 134092
rect 188956 134036 189004 134092
rect 189060 134036 189070 134092
rect 5126 133252 5136 133308
rect 5192 133252 5240 133308
rect 5296 133252 5344 133308
rect 5400 133252 5410 133308
rect 189446 133252 189456 133308
rect 189512 133252 189560 133308
rect 189616 133252 189664 133308
rect 189720 133252 189730 133308
rect 4466 132468 4476 132524
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4740 132468 4750 132524
rect 188786 132468 188796 132524
rect 188852 132468 188900 132524
rect 188956 132468 189004 132524
rect 189060 132468 189070 132524
rect 5126 131684 5136 131740
rect 5192 131684 5240 131740
rect 5296 131684 5344 131740
rect 5400 131684 5410 131740
rect 189446 131684 189456 131740
rect 189512 131684 189560 131740
rect 189616 131684 189664 131740
rect 189720 131684 189730 131740
rect 0 131348 800 131376
rect 0 131292 1708 131348
rect 1764 131292 1774 131348
rect 0 131264 800 131292
rect 4466 130900 4476 130956
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4740 130900 4750 130956
rect 188786 130900 188796 130956
rect 188852 130900 188900 130956
rect 188956 130900 189004 130956
rect 189060 130900 189070 130956
rect 5126 130116 5136 130172
rect 5192 130116 5240 130172
rect 5296 130116 5344 130172
rect 5400 130116 5410 130172
rect 189446 130116 189456 130172
rect 189512 130116 189560 130172
rect 189616 130116 189664 130172
rect 189720 130116 189730 130172
rect 4466 129332 4476 129388
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4740 129332 4750 129388
rect 188786 129332 188796 129388
rect 188852 129332 188900 129388
rect 188956 129332 189004 129388
rect 189060 129332 189070 129388
rect 5126 128548 5136 128604
rect 5192 128548 5240 128604
rect 5296 128548 5344 128604
rect 5400 128548 5410 128604
rect 189446 128548 189456 128604
rect 189512 128548 189560 128604
rect 189616 128548 189664 128604
rect 189720 128548 189730 128604
rect 205332 127988 206132 128016
rect 203746 127932 203756 127988
rect 203812 127932 206132 127988
rect 205332 127904 206132 127932
rect 4466 127764 4476 127820
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4740 127764 4750 127820
rect 188786 127764 188796 127820
rect 188852 127764 188900 127820
rect 188956 127764 189004 127820
rect 189060 127764 189070 127820
rect 0 127540 800 127568
rect 0 127484 1708 127540
rect 1764 127484 1774 127540
rect 0 127456 800 127484
rect 5126 126980 5136 127036
rect 5192 126980 5240 127036
rect 5296 126980 5344 127036
rect 5400 126980 5410 127036
rect 189446 126980 189456 127036
rect 189512 126980 189560 127036
rect 189616 126980 189664 127036
rect 189720 126980 189730 127036
rect 4466 126196 4476 126252
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4740 126196 4750 126252
rect 188786 126196 188796 126252
rect 188852 126196 188900 126252
rect 188956 126196 189004 126252
rect 189060 126196 189070 126252
rect 5126 125412 5136 125468
rect 5192 125412 5240 125468
rect 5296 125412 5344 125468
rect 5400 125412 5410 125468
rect 189446 125412 189456 125468
rect 189512 125412 189560 125468
rect 189616 125412 189664 125468
rect 189720 125412 189730 125468
rect 4466 124628 4476 124684
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4740 124628 4750 124684
rect 188786 124628 188796 124684
rect 188852 124628 188900 124684
rect 188956 124628 189004 124684
rect 189060 124628 189070 124684
rect 2818 124124 2828 124180
rect 2884 124124 26012 124180
rect 26068 124124 26078 124180
rect 5126 123844 5136 123900
rect 5192 123844 5240 123900
rect 5296 123844 5344 123900
rect 5400 123844 5410 123900
rect 189446 123844 189456 123900
rect 189512 123844 189560 123900
rect 189616 123844 189664 123900
rect 189720 123844 189730 123900
rect 0 123732 800 123760
rect 0 123676 1820 123732
rect 1876 123676 1886 123732
rect 0 123648 800 123676
rect 4466 123060 4476 123116
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4740 123060 4750 123116
rect 188786 123060 188796 123116
rect 188852 123060 188900 123116
rect 188956 123060 189004 123116
rect 189060 123060 189070 123116
rect 5126 122276 5136 122332
rect 5192 122276 5240 122332
rect 5296 122276 5344 122332
rect 5400 122276 5410 122332
rect 189446 122276 189456 122332
rect 189512 122276 189560 122332
rect 189616 122276 189664 122332
rect 189720 122276 189730 122332
rect 4466 121492 4476 121548
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4740 121492 4750 121548
rect 188786 121492 188796 121548
rect 188852 121492 188900 121548
rect 188956 121492 189004 121548
rect 189060 121492 189070 121548
rect 5126 120708 5136 120764
rect 5192 120708 5240 120764
rect 5296 120708 5344 120764
rect 5400 120708 5410 120764
rect 189446 120708 189456 120764
rect 189512 120708 189560 120764
rect 189616 120708 189664 120764
rect 189720 120708 189730 120764
rect 0 119924 800 119952
rect 4466 119924 4476 119980
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4740 119924 4750 119980
rect 188786 119924 188796 119980
rect 188852 119924 188900 119980
rect 188956 119924 189004 119980
rect 189060 119924 189070 119980
rect 0 119868 1708 119924
rect 1764 119868 1774 119924
rect 0 119840 800 119868
rect 204082 119308 204092 119364
rect 204148 119308 204260 119364
rect 204204 119252 204260 119308
rect 205332 119252 206132 119280
rect 204204 119196 206132 119252
rect 5126 119140 5136 119196
rect 5192 119140 5240 119196
rect 5296 119140 5344 119196
rect 5400 119140 5410 119196
rect 189446 119140 189456 119196
rect 189512 119140 189560 119196
rect 189616 119140 189664 119196
rect 189720 119140 189730 119196
rect 205332 119168 206132 119196
rect 202178 118636 202188 118692
rect 202244 118636 203756 118692
rect 203812 118636 203822 118692
rect 4466 118356 4476 118412
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4740 118356 4750 118412
rect 188786 118356 188796 118412
rect 188852 118356 188900 118412
rect 188956 118356 189004 118412
rect 189060 118356 189070 118412
rect 5126 117572 5136 117628
rect 5192 117572 5240 117628
rect 5296 117572 5344 117628
rect 5400 117572 5410 117628
rect 189446 117572 189456 117628
rect 189512 117572 189560 117628
rect 189616 117572 189664 117628
rect 189720 117572 189730 117628
rect 4466 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4750 116844
rect 188786 116788 188796 116844
rect 188852 116788 188900 116844
rect 188956 116788 189004 116844
rect 189060 116788 189070 116844
rect 0 116116 800 116144
rect 0 116060 1708 116116
rect 1764 116060 1774 116116
rect 0 116032 800 116060
rect 5126 116004 5136 116060
rect 5192 116004 5240 116060
rect 5296 116004 5344 116060
rect 5400 116004 5410 116060
rect 189446 116004 189456 116060
rect 189512 116004 189560 116060
rect 189616 116004 189664 116060
rect 189720 116004 189730 116060
rect 4466 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4750 115276
rect 188786 115220 188796 115276
rect 188852 115220 188900 115276
rect 188956 115220 189004 115276
rect 189060 115220 189070 115276
rect 5126 114436 5136 114492
rect 5192 114436 5240 114492
rect 5296 114436 5344 114492
rect 5400 114436 5410 114492
rect 189446 114436 189456 114492
rect 189512 114436 189560 114492
rect 189616 114436 189664 114492
rect 189720 114436 189730 114492
rect 4466 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4750 113708
rect 188786 113652 188796 113708
rect 188852 113652 188900 113708
rect 188956 113652 189004 113708
rect 189060 113652 189070 113708
rect 5126 112868 5136 112924
rect 5192 112868 5240 112924
rect 5296 112868 5344 112924
rect 5400 112868 5410 112924
rect 189446 112868 189456 112924
rect 189512 112868 189560 112924
rect 189616 112868 189664 112924
rect 189720 112868 189730 112924
rect 2818 112364 2828 112420
rect 2884 112364 9212 112420
rect 9268 112364 9278 112420
rect 0 112308 800 112336
rect 0 112252 1708 112308
rect 1764 112252 1774 112308
rect 0 112224 800 112252
rect 4466 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4750 112140
rect 188786 112084 188796 112140
rect 188852 112084 188900 112140
rect 188956 112084 189004 112140
rect 189060 112084 189070 112140
rect 5126 111300 5136 111356
rect 5192 111300 5240 111356
rect 5296 111300 5344 111356
rect 5400 111300 5410 111356
rect 189446 111300 189456 111356
rect 189512 111300 189560 111356
rect 189616 111300 189664 111356
rect 189720 111300 189730 111356
rect 4466 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4750 110572
rect 188786 110516 188796 110572
rect 188852 110516 188900 110572
rect 188956 110516 189004 110572
rect 189060 110516 189070 110572
rect 205332 110432 206132 110544
rect 5126 109732 5136 109788
rect 5192 109732 5240 109788
rect 5296 109732 5344 109788
rect 5400 109732 5410 109788
rect 189446 109732 189456 109788
rect 189512 109732 189560 109788
rect 189616 109732 189664 109788
rect 189720 109732 189730 109788
rect 4466 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4750 109004
rect 188786 108948 188796 109004
rect 188852 108948 188900 109004
rect 188956 108948 189004 109004
rect 189060 108948 189070 109004
rect 0 108500 800 108528
rect 0 108444 1708 108500
rect 1764 108444 1774 108500
rect 0 108416 800 108444
rect 5126 108164 5136 108220
rect 5192 108164 5240 108220
rect 5296 108164 5344 108220
rect 5400 108164 5410 108220
rect 189446 108164 189456 108220
rect 189512 108164 189560 108220
rect 189616 108164 189664 108220
rect 189720 108164 189730 108220
rect 4466 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4750 107436
rect 188786 107380 188796 107436
rect 188852 107380 188900 107436
rect 188956 107380 189004 107436
rect 189060 107380 189070 107436
rect 5126 106596 5136 106652
rect 5192 106596 5240 106652
rect 5296 106596 5344 106652
rect 5400 106596 5410 106652
rect 189446 106596 189456 106652
rect 189512 106596 189560 106652
rect 189616 106596 189664 106652
rect 189720 106596 189730 106652
rect 4466 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4750 105868
rect 188786 105812 188796 105868
rect 188852 105812 188900 105868
rect 188956 105812 189004 105868
rect 189060 105812 189070 105868
rect 5126 105028 5136 105084
rect 5192 105028 5240 105084
rect 5296 105028 5344 105084
rect 5400 105028 5410 105084
rect 189446 105028 189456 105084
rect 189512 105028 189560 105084
rect 189616 105028 189664 105084
rect 189720 105028 189730 105084
rect 0 104692 800 104720
rect 0 104636 1708 104692
rect 1764 104636 1774 104692
rect 0 104608 800 104636
rect 4466 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4750 104300
rect 188786 104244 188796 104300
rect 188852 104244 188900 104300
rect 188956 104244 189004 104300
rect 189060 104244 189070 104300
rect 5126 103460 5136 103516
rect 5192 103460 5240 103516
rect 5296 103460 5344 103516
rect 5400 103460 5410 103516
rect 189446 103460 189456 103516
rect 189512 103460 189560 103516
rect 189616 103460 189664 103516
rect 189720 103460 189730 103516
rect 4466 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4750 102732
rect 188786 102676 188796 102732
rect 188852 102676 188900 102732
rect 188956 102676 189004 102732
rect 189060 102676 189070 102732
rect 5126 101892 5136 101948
rect 5192 101892 5240 101948
rect 5296 101892 5344 101948
rect 5400 101892 5410 101948
rect 189446 101892 189456 101948
rect 189512 101892 189560 101948
rect 189616 101892 189664 101948
rect 189720 101892 189730 101948
rect 205332 101780 206132 101808
rect 204306 101724 204316 101780
rect 204372 101724 206132 101780
rect 205332 101696 206132 101724
rect 2034 101612 2044 101668
rect 2100 101612 7532 101668
rect 7588 101612 7598 101668
rect 1698 101388 1708 101444
rect 1764 101388 2492 101444
rect 2548 101388 2558 101444
rect 4466 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4750 101164
rect 188786 101108 188796 101164
rect 188852 101108 188900 101164
rect 188956 101108 189004 101164
rect 189060 101108 189070 101164
rect 0 100884 800 100912
rect 0 100828 1708 100884
rect 1764 100828 1774 100884
rect 0 100800 800 100828
rect 5126 100324 5136 100380
rect 5192 100324 5240 100380
rect 5296 100324 5344 100380
rect 5400 100324 5410 100380
rect 189446 100324 189456 100380
rect 189512 100324 189560 100380
rect 189616 100324 189664 100380
rect 189720 100324 189730 100380
rect 4466 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4750 99596
rect 188786 99540 188796 99596
rect 188852 99540 188900 99596
rect 188956 99540 189004 99596
rect 189060 99540 189070 99596
rect 5126 98756 5136 98812
rect 5192 98756 5240 98812
rect 5296 98756 5344 98812
rect 5400 98756 5410 98812
rect 189446 98756 189456 98812
rect 189512 98756 189560 98812
rect 189616 98756 189664 98812
rect 189720 98756 189730 98812
rect 4466 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4750 98028
rect 188786 97972 188796 98028
rect 188852 97972 188900 98028
rect 188956 97972 189004 98028
rect 189060 97972 189070 98028
rect 5126 97188 5136 97244
rect 5192 97188 5240 97244
rect 5296 97188 5344 97244
rect 5400 97188 5410 97244
rect 189446 97188 189456 97244
rect 189512 97188 189560 97244
rect 189616 97188 189664 97244
rect 189720 97188 189730 97244
rect 0 97076 800 97104
rect 0 97020 1708 97076
rect 1764 97020 1774 97076
rect 0 96992 800 97020
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 188786 96404 188796 96460
rect 188852 96404 188900 96460
rect 188956 96404 189004 96460
rect 189060 96404 189070 96460
rect 5126 95620 5136 95676
rect 5192 95620 5240 95676
rect 5296 95620 5344 95676
rect 5400 95620 5410 95676
rect 189446 95620 189456 95676
rect 189512 95620 189560 95676
rect 189616 95620 189664 95676
rect 189720 95620 189730 95676
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 188786 94836 188796 94892
rect 188852 94836 188900 94892
rect 188956 94836 189004 94892
rect 189060 94836 189070 94892
rect 5126 94052 5136 94108
rect 5192 94052 5240 94108
rect 5296 94052 5344 94108
rect 5400 94052 5410 94108
rect 189446 94052 189456 94108
rect 189512 94052 189560 94108
rect 189616 94052 189664 94108
rect 189720 94052 189730 94108
rect 190642 93660 190652 93716
rect 190708 93660 201180 93716
rect 201236 93660 203980 93716
rect 204036 93660 204046 93716
rect 1698 93436 1708 93492
rect 1764 93436 1774 93492
rect 0 93268 800 93296
rect 1708 93268 1764 93436
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 188786 93268 188796 93324
rect 188852 93268 188900 93324
rect 188956 93268 189004 93324
rect 189060 93268 189070 93324
rect 0 93212 1764 93268
rect 0 93184 800 93212
rect 205332 93044 206132 93072
rect 203186 92988 203196 93044
rect 203252 92988 206132 93044
rect 205332 92960 206132 92988
rect 5126 92484 5136 92540
rect 5192 92484 5240 92540
rect 5296 92484 5344 92540
rect 5400 92484 5410 92540
rect 189446 92484 189456 92540
rect 189512 92484 189560 92540
rect 189616 92484 189664 92540
rect 189720 92484 189730 92540
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 188786 91700 188796 91756
rect 188852 91700 188900 91756
rect 188956 91700 189004 91756
rect 189060 91700 189070 91756
rect 5126 90916 5136 90972
rect 5192 90916 5240 90972
rect 5296 90916 5344 90972
rect 5400 90916 5410 90972
rect 189446 90916 189456 90972
rect 189512 90916 189560 90972
rect 189616 90916 189664 90972
rect 189720 90916 189730 90972
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 188786 90132 188796 90188
rect 188852 90132 188900 90188
rect 188956 90132 189004 90188
rect 189060 90132 189070 90188
rect 0 89460 800 89488
rect 0 89404 1708 89460
rect 1764 89404 2492 89460
rect 2548 89404 2558 89460
rect 0 89376 800 89404
rect 5126 89348 5136 89404
rect 5192 89348 5240 89404
rect 5296 89348 5344 89404
rect 5400 89348 5410 89404
rect 189446 89348 189456 89404
rect 189512 89348 189560 89404
rect 189616 89348 189664 89404
rect 189720 89348 189730 89404
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 188786 88564 188796 88620
rect 188852 88564 188900 88620
rect 188956 88564 189004 88620
rect 189060 88564 189070 88620
rect 5126 87780 5136 87836
rect 5192 87780 5240 87836
rect 5296 87780 5344 87836
rect 5400 87780 5410 87836
rect 189446 87780 189456 87836
rect 189512 87780 189560 87836
rect 189616 87780 189664 87836
rect 189720 87780 189730 87836
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 188786 86996 188796 87052
rect 188852 86996 188900 87052
rect 188956 86996 189004 87052
rect 189060 86996 189070 87052
rect 5126 86212 5136 86268
rect 5192 86212 5240 86268
rect 5296 86212 5344 86268
rect 5400 86212 5410 86268
rect 189446 86212 189456 86268
rect 189512 86212 189560 86268
rect 189616 86212 189664 86268
rect 189720 86212 189730 86268
rect 0 85652 800 85680
rect 0 85596 1708 85652
rect 1764 85596 1774 85652
rect 0 85568 800 85596
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 188786 85428 188796 85484
rect 188852 85428 188900 85484
rect 188956 85428 189004 85484
rect 189060 85428 189070 85484
rect 5126 84644 5136 84700
rect 5192 84644 5240 84700
rect 5296 84644 5344 84700
rect 5400 84644 5410 84700
rect 189446 84644 189456 84700
rect 189512 84644 189560 84700
rect 189616 84644 189664 84700
rect 189720 84644 189730 84700
rect 205332 84224 206132 84336
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 188786 83860 188796 83916
rect 188852 83860 188900 83916
rect 188956 83860 189004 83916
rect 189060 83860 189070 83916
rect 5126 83076 5136 83132
rect 5192 83076 5240 83132
rect 5296 83076 5344 83132
rect 5400 83076 5410 83132
rect 189446 83076 189456 83132
rect 189512 83076 189560 83132
rect 189616 83076 189664 83132
rect 189720 83076 189730 83132
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 188786 82292 188796 82348
rect 188852 82292 188900 82348
rect 188956 82292 189004 82348
rect 189060 82292 189070 82348
rect 1698 82012 1708 82068
rect 1764 82012 1774 82068
rect 0 81844 800 81872
rect 1708 81844 1764 82012
rect 0 81788 1764 81844
rect 0 81760 800 81788
rect 5126 81508 5136 81564
rect 5192 81508 5240 81564
rect 5296 81508 5344 81564
rect 5400 81508 5410 81564
rect 189446 81508 189456 81564
rect 189512 81508 189560 81564
rect 189616 81508 189664 81564
rect 189720 81508 189730 81564
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 188786 80724 188796 80780
rect 188852 80724 188900 80780
rect 188956 80724 189004 80780
rect 189060 80724 189070 80780
rect 5126 79940 5136 79996
rect 5192 79940 5240 79996
rect 5296 79940 5344 79996
rect 5400 79940 5410 79996
rect 189446 79940 189456 79996
rect 189512 79940 189560 79996
rect 189616 79940 189664 79996
rect 189720 79940 189730 79996
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 188786 79156 188796 79212
rect 188852 79156 188900 79212
rect 188956 79156 189004 79212
rect 189060 79156 189070 79212
rect 1698 78540 1708 78596
rect 1764 78540 2492 78596
rect 2548 78540 2558 78596
rect 14242 78540 14252 78596
rect 14308 78540 17612 78596
rect 17668 78540 20132 78596
rect 5126 78372 5136 78428
rect 5192 78372 5240 78428
rect 5296 78372 5344 78428
rect 5400 78372 5410 78428
rect 20076 78382 20132 78540
rect 189446 78372 189456 78428
rect 189512 78372 189560 78428
rect 189616 78372 189664 78428
rect 189720 78372 189730 78428
rect 0 78036 800 78064
rect 0 77980 1708 78036
rect 1764 77980 1774 78036
rect 0 77952 800 77980
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 188786 77588 188796 77644
rect 188852 77588 188900 77644
rect 188956 77588 189004 77644
rect 189060 77588 189070 77644
rect 5126 76804 5136 76860
rect 5192 76804 5240 76860
rect 5296 76804 5344 76860
rect 5400 76804 5410 76860
rect 20076 76580 20132 77194
rect 189446 76804 189456 76860
rect 189512 76804 189560 76860
rect 189616 76804 189664 76860
rect 189720 76804 189730 76860
rect 15922 76524 15932 76580
rect 15988 76524 17612 76580
rect 17668 76524 20132 76580
rect 2258 76300 2268 76356
rect 2324 76300 17612 76356
rect 17668 76300 20132 76356
rect 20076 76270 20132 76300
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 188786 76020 188796 76076
rect 188852 76020 188900 76076
rect 188956 76020 189004 76076
rect 189060 76020 189070 76076
rect 2034 75628 2044 75684
rect 2100 75628 17500 75684
rect 17556 75628 20244 75684
rect 5126 75236 5136 75292
rect 5192 75236 5240 75292
rect 5296 75236 5344 75292
rect 5400 75236 5410 75292
rect 20188 75082 20244 75628
rect 205332 75572 206132 75600
rect 204306 75516 204316 75572
rect 204372 75516 206132 75572
rect 205332 75488 206132 75516
rect 189446 75236 189456 75292
rect 189512 75236 189560 75292
rect 189616 75236 189664 75292
rect 189720 75236 189730 75292
rect 2146 74732 2156 74788
rect 2212 74732 17500 74788
rect 17556 74732 20132 74788
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 20076 74290 20132 74732
rect 188786 74452 188796 74508
rect 188852 74452 188900 74508
rect 188956 74452 189004 74508
rect 189060 74452 189070 74508
rect 0 74228 800 74256
rect 0 74172 1708 74228
rect 1764 74172 1774 74228
rect 0 74144 800 74172
rect 5126 73668 5136 73724
rect 5192 73668 5240 73724
rect 5296 73668 5344 73724
rect 5400 73668 5410 73724
rect 189446 73668 189456 73724
rect 189512 73668 189560 73724
rect 189616 73668 189664 73724
rect 189720 73668 189730 73724
rect 20076 73220 20132 73234
rect 7522 73164 7532 73220
rect 7588 73164 17500 73220
rect 17556 73164 20132 73220
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 188786 72884 188796 72940
rect 188852 72884 188900 72940
rect 188956 72884 189004 72940
rect 189060 72884 189070 72940
rect 5126 72100 5136 72156
rect 5192 72100 5240 72156
rect 5296 72100 5344 72156
rect 5400 72100 5410 72156
rect 189446 72100 189456 72156
rect 189512 72100 189560 72156
rect 189616 72100 189664 72156
rect 189720 72100 189730 72156
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 188786 71316 188796 71372
rect 188852 71316 188900 71372
rect 188956 71316 189004 71372
rect 189060 71316 189070 71372
rect 5126 70532 5136 70588
rect 5192 70532 5240 70588
rect 5296 70532 5344 70588
rect 5400 70532 5410 70588
rect 189446 70532 189456 70588
rect 189512 70532 189560 70588
rect 189616 70532 189664 70588
rect 189720 70532 189730 70588
rect 0 70420 800 70448
rect 0 70364 1708 70420
rect 1764 70364 1774 70420
rect 0 70336 800 70364
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 188786 69748 188796 69804
rect 188852 69748 188900 69804
rect 188956 69748 189004 69804
rect 189060 69748 189070 69804
rect 5126 68964 5136 69020
rect 5192 68964 5240 69020
rect 5296 68964 5344 69020
rect 5400 68964 5410 69020
rect 189446 68964 189456 69020
rect 189512 68964 189560 69020
rect 189616 68964 189664 69020
rect 189720 68964 189730 69020
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 188786 68180 188796 68236
rect 188852 68180 188900 68236
rect 188956 68180 189004 68236
rect 189060 68180 189070 68236
rect 5126 67396 5136 67452
rect 5192 67396 5240 67452
rect 5296 67396 5344 67452
rect 5400 67396 5410 67452
rect 189446 67396 189456 67452
rect 189512 67396 189560 67452
rect 189616 67396 189664 67452
rect 189720 67396 189730 67452
rect 187282 67004 187292 67060
rect 187348 67004 201180 67060
rect 201236 67004 203980 67060
rect 204036 67004 204046 67060
rect 205332 66836 206132 66864
rect 203186 66780 203196 66836
rect 203252 66780 206132 66836
rect 205332 66752 206132 66780
rect 0 66612 800 66640
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 188786 66612 188796 66668
rect 188852 66612 188900 66668
rect 188956 66612 189004 66668
rect 189060 66612 189070 66668
rect 0 66556 1708 66612
rect 1764 66556 2492 66612
rect 2548 66556 2558 66612
rect 0 66528 800 66556
rect 5126 65828 5136 65884
rect 5192 65828 5240 65884
rect 5296 65828 5344 65884
rect 5400 65828 5410 65884
rect 189446 65828 189456 65884
rect 189512 65828 189560 65884
rect 189616 65828 189664 65884
rect 189720 65828 189730 65884
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 188786 65044 188796 65100
rect 188852 65044 188900 65100
rect 188956 65044 189004 65100
rect 189060 65044 189070 65100
rect 5126 64260 5136 64316
rect 5192 64260 5240 64316
rect 5296 64260 5344 64316
rect 5400 64260 5410 64316
rect 189446 64260 189456 64316
rect 189512 64260 189560 64316
rect 189616 64260 189664 64316
rect 189720 64260 189730 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 188786 63476 188796 63532
rect 188852 63476 188900 63532
rect 188956 63476 189004 63532
rect 189060 63476 189070 63532
rect 1698 62860 1708 62916
rect 1764 62860 1774 62916
rect 0 62804 800 62832
rect 1708 62804 1764 62860
rect 0 62748 1764 62804
rect 0 62720 800 62748
rect 5126 62692 5136 62748
rect 5192 62692 5240 62748
rect 5296 62692 5344 62748
rect 5400 62692 5410 62748
rect 189446 62692 189456 62748
rect 189512 62692 189560 62748
rect 189616 62692 189664 62748
rect 189720 62692 189730 62748
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 188786 61908 188796 61964
rect 188852 61908 188900 61964
rect 188956 61908 189004 61964
rect 189060 61908 189070 61964
rect 5126 61124 5136 61180
rect 5192 61124 5240 61180
rect 5296 61124 5344 61180
rect 5400 61124 5410 61180
rect 189446 61124 189456 61180
rect 189512 61124 189560 61180
rect 189616 61124 189664 61180
rect 189720 61124 189730 61180
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 188786 60340 188796 60396
rect 188852 60340 188900 60396
rect 188956 60340 189004 60396
rect 189060 60340 189070 60396
rect 5126 59556 5136 59612
rect 5192 59556 5240 59612
rect 5296 59556 5344 59612
rect 5400 59556 5410 59612
rect 189446 59556 189456 59612
rect 189512 59556 189560 59612
rect 189616 59556 189664 59612
rect 189720 59556 189730 59612
rect 0 58996 800 59024
rect 0 58940 1708 58996
rect 1764 58940 1774 58996
rect 0 58912 800 58940
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 188786 58772 188796 58828
rect 188852 58772 188900 58828
rect 188956 58772 189004 58828
rect 189060 58772 189070 58828
rect 5126 57988 5136 58044
rect 5192 57988 5240 58044
rect 5296 57988 5344 58044
rect 5400 57988 5410 58044
rect 189446 57988 189456 58044
rect 189512 57988 189560 58044
rect 189616 57988 189664 58044
rect 189720 57988 189730 58044
rect 205332 58016 206132 58128
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 188786 57204 188796 57260
rect 188852 57204 188900 57260
rect 188956 57204 189004 57260
rect 189060 57204 189070 57260
rect 5126 56420 5136 56476
rect 5192 56420 5240 56476
rect 5296 56420 5344 56476
rect 5400 56420 5410 56476
rect 189446 56420 189456 56476
rect 189512 56420 189560 56476
rect 189616 56420 189664 56476
rect 189720 56420 189730 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 188786 55636 188796 55692
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 189060 55636 189070 55692
rect 2258 55244 2268 55300
rect 2324 55244 15932 55300
rect 15988 55244 15998 55300
rect 0 55188 800 55216
rect 0 55132 1708 55188
rect 1764 55132 1774 55188
rect 0 55104 800 55132
rect 5126 54852 5136 54908
rect 5192 54852 5240 54908
rect 5296 54852 5344 54908
rect 5400 54852 5410 54908
rect 189446 54852 189456 54908
rect 189512 54852 189560 54908
rect 189616 54852 189664 54908
rect 189720 54852 189730 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 188786 54068 188796 54124
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 189060 54068 189070 54124
rect 5126 53284 5136 53340
rect 5192 53284 5240 53340
rect 5296 53284 5344 53340
rect 5400 53284 5410 53340
rect 189446 53284 189456 53340
rect 189512 53284 189560 53340
rect 189616 53284 189664 53340
rect 189720 53284 189730 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 188786 52500 188796 52556
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 189060 52500 189070 52556
rect 5126 51716 5136 51772
rect 5192 51716 5240 51772
rect 5296 51716 5344 51772
rect 5400 51716 5410 51772
rect 189446 51716 189456 51772
rect 189512 51716 189560 51772
rect 189616 51716 189664 51772
rect 189720 51716 189730 51772
rect 0 51380 800 51408
rect 0 51324 1708 51380
rect 1764 51324 1774 51380
rect 0 51296 800 51324
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 188786 50932 188796 50988
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 189060 50932 189070 50988
rect 5126 50148 5136 50204
rect 5192 50148 5240 50204
rect 5296 50148 5344 50204
rect 5400 50148 5410 50204
rect 189446 50148 189456 50204
rect 189512 50148 189560 50204
rect 189616 50148 189664 50204
rect 189720 50148 189730 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 188786 49364 188796 49420
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 189060 49364 189070 49420
rect 205332 49364 206132 49392
rect 203746 49308 203756 49364
rect 203812 49308 206132 49364
rect 205332 49280 206132 49308
rect 5126 48580 5136 48636
rect 5192 48580 5240 48636
rect 5296 48580 5344 48636
rect 5400 48580 5410 48636
rect 189446 48580 189456 48636
rect 189512 48580 189560 48636
rect 189616 48580 189664 48636
rect 189720 48580 189730 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 188786 47796 188796 47852
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 189060 47796 189070 47852
rect 0 47572 800 47600
rect 0 47516 1708 47572
rect 1764 47516 1774 47572
rect 0 47488 800 47516
rect 5126 47012 5136 47068
rect 5192 47012 5240 47068
rect 5296 47012 5344 47068
rect 5400 47012 5410 47068
rect 189446 47012 189456 47068
rect 189512 47012 189560 47068
rect 189616 47012 189664 47068
rect 189720 47012 189730 47068
rect 132934 46956 132972 47012
rect 133028 46956 133038 47012
rect 156342 46956 156380 47012
rect 156436 46956 156446 47012
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 188786 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189070 46284
rect 132934 45724 132972 45780
rect 133028 45724 133038 45780
rect 156342 45724 156380 45780
rect 156436 45724 156446 45780
rect 5126 45444 5136 45500
rect 5192 45444 5240 45500
rect 5296 45444 5344 45500
rect 5400 45444 5410 45500
rect 189446 45444 189456 45500
rect 189512 45444 189560 45500
rect 189616 45444 189664 45500
rect 189720 45444 189730 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 188786 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189070 44716
rect 2258 44268 2268 44324
rect 2324 44268 14252 44324
rect 14308 44268 14318 44324
rect 5126 43876 5136 43932
rect 5192 43876 5240 43932
rect 5296 43876 5344 43932
rect 5400 43876 5410 43932
rect 189446 43876 189456 43932
rect 189512 43876 189560 43932
rect 189616 43876 189664 43932
rect 189720 43876 189730 43932
rect 0 43764 800 43792
rect 0 43708 1820 43764
rect 1876 43708 1886 43764
rect 0 43680 800 43708
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 188786 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189070 43148
rect 5126 42308 5136 42364
rect 5192 42308 5240 42364
rect 5296 42308 5344 42364
rect 5400 42308 5410 42364
rect 189446 42308 189456 42364
rect 189512 42308 189560 42364
rect 189616 42308 189664 42364
rect 189720 42308 189730 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 188786 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189070 41580
rect 64418 41244 64428 41300
rect 64484 41244 71932 41300
rect 71988 41244 71998 41300
rect 56242 41132 56252 41188
rect 56308 41132 75516 41188
rect 75572 41132 75582 41188
rect 63746 41020 63756 41076
rect 63812 41020 67676 41076
rect 67732 41020 67742 41076
rect 85138 40908 85148 40964
rect 85204 40908 201404 40964
rect 201460 40908 201470 40964
rect 5126 40740 5136 40796
rect 5192 40740 5240 40796
rect 5296 40740 5344 40796
rect 5400 40740 5410 40796
rect 189446 40740 189456 40796
rect 189512 40740 189560 40796
rect 189616 40740 189664 40796
rect 189720 40740 189730 40796
rect 205332 40628 206132 40656
rect 204082 40572 204092 40628
rect 204148 40572 206132 40628
rect 205332 40544 206132 40572
rect 0 39956 800 39984
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 188786 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189070 40012
rect 0 39900 1708 39956
rect 1764 39900 1774 39956
rect 0 39872 800 39900
rect 5126 39172 5136 39228
rect 5192 39172 5240 39228
rect 5296 39172 5344 39228
rect 5400 39172 5410 39228
rect 189446 39172 189456 39228
rect 189512 39172 189560 39228
rect 189616 39172 189664 39228
rect 189720 39172 189730 39228
rect 173954 38668 173964 38724
rect 174020 38668 188748 38724
rect 188804 38668 188814 38724
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 61730 38108 61740 38164
rect 61796 38108 132972 38164
rect 133028 38108 133038 38164
rect 26002 37996 26012 38052
rect 26068 37996 51436 38052
rect 51492 37996 51502 38052
rect 59042 37996 59052 38052
rect 59108 37996 156380 38052
rect 156436 37996 156446 38052
rect 184716 37726 184772 38668
rect 188786 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189070 38444
rect 5126 37604 5136 37660
rect 5192 37604 5240 37660
rect 5296 37604 5344 37660
rect 5400 37604 5410 37660
rect 189446 37604 189456 37660
rect 189512 37604 189560 37660
rect 189616 37604 189664 37660
rect 189720 37604 189730 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 188786 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189070 36876
rect 20076 36260 20132 36274
rect 2034 36204 2044 36260
rect 2100 36204 17612 36260
rect 17668 36204 20132 36260
rect 0 36148 800 36176
rect 0 36092 1708 36148
rect 1764 36092 1774 36148
rect 0 36064 800 36092
rect 5126 36036 5136 36092
rect 5192 36036 5240 36092
rect 5296 36036 5344 36092
rect 5400 36036 5410 36092
rect 189446 36036 189456 36092
rect 189512 36036 189560 36092
rect 189616 36036 189664 36092
rect 189720 36036 189730 36092
rect 12674 35532 12684 35588
rect 12740 35532 17612 35588
rect 17668 35532 19460 35588
rect 19404 35510 19460 35532
rect 19404 35454 20104 35510
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 188786 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189070 35308
rect 20076 34692 20132 35218
rect 2146 34636 2156 34692
rect 2212 34636 16940 34692
rect 16996 34636 20132 34692
rect 5126 34468 5136 34524
rect 5192 34468 5240 34524
rect 5296 34468 5344 34524
rect 5400 34468 5410 34524
rect 189446 34468 189456 34524
rect 189512 34468 189560 34524
rect 189616 34468 189664 34524
rect 189720 34468 189730 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 188786 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189070 33740
rect 5126 32900 5136 32956
rect 5192 32900 5240 32956
rect 5296 32900 5344 32956
rect 5400 32900 5410 32956
rect 189446 32900 189456 32956
rect 189512 32900 189560 32956
rect 189616 32900 189664 32956
rect 189720 32900 189730 32956
rect 0 32340 800 32368
rect 0 32284 1708 32340
rect 1764 32284 2492 32340
rect 2548 32284 2558 32340
rect 0 32256 800 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 188786 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189070 32172
rect 82338 31836 82348 31892
rect 82404 31836 85148 31892
rect 85204 31836 85214 31892
rect 205332 31808 206132 31920
rect 5126 31332 5136 31388
rect 5192 31332 5240 31388
rect 5296 31332 5344 31388
rect 5400 31332 5410 31388
rect 189446 31332 189456 31388
rect 189512 31332 189560 31388
rect 189616 31332 189664 31388
rect 189720 31332 189730 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 188786 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189070 30604
rect 5126 29764 5136 29820
rect 5192 29764 5240 29820
rect 5296 29764 5344 29820
rect 5400 29764 5410 29820
rect 189446 29764 189456 29820
rect 189512 29764 189560 29820
rect 189616 29764 189664 29820
rect 189720 29764 189730 29820
rect 2370 29372 2380 29428
rect 2436 29372 75628 29428
rect 75684 29372 75694 29428
rect 154578 29372 154588 29428
rect 154644 29372 196588 29428
rect 196644 29372 196654 29428
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 188786 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189070 29036
rect 0 28532 800 28560
rect 0 28476 1708 28532
rect 1764 28476 1774 28532
rect 0 28448 800 28476
rect 5126 28196 5136 28252
rect 5192 28196 5240 28252
rect 5296 28196 5344 28252
rect 5400 28196 5410 28252
rect 189446 28196 189456 28252
rect 189512 28196 189560 28252
rect 189616 28196 189664 28252
rect 189720 28196 189730 28252
rect 154690 27804 154700 27860
rect 154756 27804 201068 27860
rect 201124 27804 201134 27860
rect 9202 27692 9212 27748
rect 9268 27692 53900 27748
rect 53956 27692 53966 27748
rect 155138 27692 155148 27748
rect 155204 27692 202412 27748
rect 202468 27692 202478 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 188786 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189070 27468
rect 5126 26628 5136 26684
rect 5192 26628 5240 26684
rect 5296 26628 5344 26684
rect 5400 26628 5410 26684
rect 189446 26628 189456 26684
rect 189512 26628 189560 26684
rect 189616 26628 189664 26684
rect 189720 26628 189730 26684
rect 140018 26124 140028 26180
rect 140084 26124 149548 26180
rect 149604 26124 154700 26180
rect 154756 26124 154766 26180
rect 125346 26012 125356 26068
rect 125412 26012 154812 26068
rect 154868 26012 155148 26068
rect 155204 26012 155214 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 188786 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189070 25900
rect 102452 25564 187292 25620
rect 187348 25564 187358 25620
rect 102452 25508 102508 25564
rect 78866 25452 78876 25508
rect 78932 25452 96572 25508
rect 96628 25452 102508 25508
rect 77186 25340 77196 25396
rect 77252 25340 110908 25396
rect 110964 25340 190652 25396
rect 190708 25340 190718 25396
rect 78642 25228 78652 25284
rect 78708 25228 82012 25284
rect 82068 25228 82078 25284
rect 5126 25060 5136 25116
rect 5192 25060 5240 25116
rect 5296 25060 5344 25116
rect 5400 25060 5410 25116
rect 189446 25060 189456 25116
rect 189512 25060 189560 25116
rect 189616 25060 189664 25116
rect 189720 25060 189730 25116
rect 0 24724 800 24752
rect 0 24668 1708 24724
rect 1764 24668 1774 24724
rect 0 24640 800 24668
rect 12562 24332 12572 24388
rect 12628 24332 44156 24388
rect 44212 24332 44222 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 188786 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189070 24332
rect 5126 23492 5136 23548
rect 5192 23492 5240 23548
rect 5296 23492 5344 23548
rect 5400 23492 5410 23548
rect 189446 23492 189456 23548
rect 189512 23492 189560 23548
rect 189616 23492 189664 23548
rect 189720 23492 189730 23548
rect 205332 23156 206132 23184
rect 204306 23100 204316 23156
rect 204372 23100 206132 23156
rect 205332 23072 206132 23100
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 149492 22708 149548 22932
rect 149604 22876 149614 22932
rect 188786 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189070 22764
rect 78866 22652 78876 22708
rect 78932 22652 97132 22708
rect 97188 22652 97198 22708
rect 140018 22652 140028 22708
rect 140084 22652 149548 22708
rect 51426 22316 51436 22372
rect 51492 22316 51502 22372
rect 61730 22316 61740 22372
rect 61796 22316 61806 22372
rect 65090 22316 65100 22372
rect 65156 22316 65268 22372
rect 71922 22316 71932 22372
rect 71988 22316 72100 22372
rect 51436 22120 51492 22316
rect 61740 22120 61796 22316
rect 65212 22120 65268 22316
rect 72044 22120 72100 22316
rect 5126 21924 5136 21980
rect 5192 21924 5240 21980
rect 5296 21924 5344 21980
rect 5400 21924 5410 21980
rect 189446 21924 189456 21980
rect 189512 21924 189560 21980
rect 189616 21924 189664 21980
rect 189720 21924 189730 21980
rect 44118 21756 44156 21812
rect 44212 21756 44222 21812
rect 53890 21756 53900 21812
rect 53956 21756 54348 21812
rect 54404 21756 54414 21812
rect 67666 21756 67676 21812
rect 67732 21756 68348 21812
rect 68404 21756 68796 21812
rect 68852 21756 68862 21812
rect 75282 21756 75292 21812
rect 75348 21756 75516 21812
rect 75572 21756 75582 21812
rect 55094 21644 55132 21700
rect 55188 21644 55198 21700
rect 1698 21420 1708 21476
rect 1764 21420 2492 21476
rect 2548 21420 2558 21476
rect 44678 21196 44716 21252
rect 44772 21196 44782 21252
rect 78642 21196 78652 21252
rect 78708 21196 82908 21252
rect 82964 21196 82974 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 188786 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189070 21196
rect 77186 21084 77196 21140
rect 77252 21084 111244 21140
rect 111300 21084 111310 21140
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 0 20832 800 20860
rect 17714 20412 17724 20468
rect 17780 20412 48300 20468
rect 48356 20412 48366 20468
rect 67750 20412 67788 20468
rect 67844 20412 67854 20468
rect 75618 20412 75628 20468
rect 75684 20412 82460 20468
rect 82516 20412 82526 20468
rect 154242 20412 154252 20468
rect 154308 20412 154588 20468
rect 154644 20412 154654 20468
rect 5126 20356 5136 20412
rect 5192 20356 5240 20412
rect 5296 20356 5344 20412
rect 5400 20356 5410 20412
rect 189446 20356 189456 20412
rect 189512 20356 189560 20412
rect 189616 20356 189664 20412
rect 189720 20356 189730 20412
rect 58706 19852 58716 19908
rect 58772 19852 59052 19908
rect 59108 19852 59118 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 188786 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189070 19628
rect 5126 18788 5136 18844
rect 5192 18788 5240 18844
rect 5296 18788 5344 18844
rect 5400 18788 5410 18844
rect 189446 18788 189456 18844
rect 189512 18788 189560 18844
rect 189616 18788 189664 18844
rect 189720 18788 189730 18844
rect 22754 18396 22764 18452
rect 22820 18396 77308 18452
rect 77364 18396 77374 18452
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 188786 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189070 18060
rect 5126 17220 5136 17276
rect 5192 17220 5240 17276
rect 5296 17220 5344 17276
rect 5400 17220 5410 17276
rect 35846 17220 35856 17276
rect 35912 17220 35960 17276
rect 36016 17220 36064 17276
rect 36120 17220 36130 17276
rect 66566 17220 66576 17276
rect 66632 17220 66680 17276
rect 66736 17220 66784 17276
rect 66840 17220 66850 17276
rect 97286 17220 97296 17276
rect 97352 17220 97400 17276
rect 97456 17220 97504 17276
rect 97560 17220 97570 17276
rect 128006 17220 128016 17276
rect 128072 17220 128120 17276
rect 128176 17220 128224 17276
rect 128280 17220 128290 17276
rect 158726 17220 158736 17276
rect 158792 17220 158840 17276
rect 158896 17220 158944 17276
rect 159000 17220 159010 17276
rect 189446 17220 189456 17276
rect 189512 17220 189560 17276
rect 189616 17220 189664 17276
rect 189720 17220 189730 17276
rect 0 17108 800 17136
rect 0 17052 1708 17108
rect 1764 17052 1774 17108
rect 77298 17052 77308 17108
rect 77364 17052 78876 17108
rect 78932 17052 78988 17108
rect 79044 17052 79054 17108
rect 0 17024 800 17052
rect 125570 16828 125580 16884
rect 125636 16828 154812 16884
rect 154868 16828 154878 16884
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 127346 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127630 16492
rect 158066 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158350 16492
rect 188786 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189070 16492
rect 5126 15652 5136 15708
rect 5192 15652 5240 15708
rect 5296 15652 5344 15708
rect 5400 15652 5410 15708
rect 35846 15652 35856 15708
rect 35912 15652 35960 15708
rect 36016 15652 36064 15708
rect 36120 15652 36130 15708
rect 66566 15652 66576 15708
rect 66632 15652 66680 15708
rect 66736 15652 66784 15708
rect 66840 15652 66850 15708
rect 97286 15652 97296 15708
rect 97352 15652 97400 15708
rect 97456 15652 97504 15708
rect 97560 15652 97570 15708
rect 128006 15652 128016 15708
rect 128072 15652 128120 15708
rect 128176 15652 128224 15708
rect 128280 15652 128290 15708
rect 158726 15652 158736 15708
rect 158792 15652 158840 15708
rect 158896 15652 158944 15708
rect 159000 15652 159010 15708
rect 189446 15652 189456 15708
rect 189512 15652 189560 15708
rect 189616 15652 189664 15708
rect 189720 15652 189730 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 127346 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127630 14924
rect 158066 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158350 14924
rect 188786 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189070 14924
rect 67890 14476 67900 14532
rect 67956 14476 201740 14532
rect 201796 14476 204316 14532
rect 204372 14476 204382 14532
rect 205332 14420 206132 14448
rect 204082 14364 204092 14420
rect 204148 14364 206132 14420
rect 205332 14336 206132 14364
rect 5126 14084 5136 14140
rect 5192 14084 5240 14140
rect 5296 14084 5344 14140
rect 5400 14084 5410 14140
rect 35846 14084 35856 14140
rect 35912 14084 35960 14140
rect 36016 14084 36064 14140
rect 36120 14084 36130 14140
rect 66566 14084 66576 14140
rect 66632 14084 66680 14140
rect 66736 14084 66784 14140
rect 66840 14084 66850 14140
rect 97286 14084 97296 14140
rect 97352 14084 97400 14140
rect 97456 14084 97504 14140
rect 97560 14084 97570 14140
rect 128006 14084 128016 14140
rect 128072 14084 128120 14140
rect 128176 14084 128224 14140
rect 128280 14084 128290 14140
rect 158726 14084 158736 14140
rect 158792 14084 158840 14140
rect 158896 14084 158944 14140
rect 159000 14084 159010 14140
rect 189446 14084 189456 14140
rect 189512 14084 189560 14140
rect 189616 14084 189664 14140
rect 189720 14084 189730 14140
rect 0 13300 800 13328
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 127346 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127630 13356
rect 158066 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158350 13356
rect 188786 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189070 13356
rect 0 13244 1708 13300
rect 1764 13244 1774 13300
rect 0 13216 800 13244
rect 5126 12516 5136 12572
rect 5192 12516 5240 12572
rect 5296 12516 5344 12572
rect 5400 12516 5410 12572
rect 35846 12516 35856 12572
rect 35912 12516 35960 12572
rect 36016 12516 36064 12572
rect 36120 12516 36130 12572
rect 66566 12516 66576 12572
rect 66632 12516 66680 12572
rect 66736 12516 66784 12572
rect 66840 12516 66850 12572
rect 97286 12516 97296 12572
rect 97352 12516 97400 12572
rect 97456 12516 97504 12572
rect 97560 12516 97570 12572
rect 128006 12516 128016 12572
rect 128072 12516 128120 12572
rect 128176 12516 128224 12572
rect 128280 12516 128290 12572
rect 158726 12516 158736 12572
rect 158792 12516 158840 12572
rect 158896 12516 158944 12572
rect 159000 12516 159010 12572
rect 189446 12516 189456 12572
rect 189512 12516 189560 12572
rect 189616 12516 189664 12572
rect 189720 12516 189730 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 127346 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127630 11788
rect 158066 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158350 11788
rect 188786 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189070 11788
rect 5126 10948 5136 11004
rect 5192 10948 5240 11004
rect 5296 10948 5344 11004
rect 5400 10948 5410 11004
rect 35846 10948 35856 11004
rect 35912 10948 35960 11004
rect 36016 10948 36064 11004
rect 36120 10948 36130 11004
rect 66566 10948 66576 11004
rect 66632 10948 66680 11004
rect 66736 10948 66784 11004
rect 66840 10948 66850 11004
rect 97286 10948 97296 11004
rect 97352 10948 97400 11004
rect 97456 10948 97504 11004
rect 97560 10948 97570 11004
rect 128006 10948 128016 11004
rect 128072 10948 128120 11004
rect 128176 10948 128224 11004
rect 128280 10948 128290 11004
rect 158726 10948 158736 11004
rect 158792 10948 158840 11004
rect 158896 10948 158944 11004
rect 159000 10948 159010 11004
rect 189446 10948 189456 11004
rect 189512 10948 189560 11004
rect 189616 10948 189664 11004
rect 189720 10948 189730 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 127346 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127630 10220
rect 158066 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158350 10220
rect 188786 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189070 10220
rect 2034 9548 2044 9604
rect 2100 9548 12684 9604
rect 12740 9548 12750 9604
rect 0 9492 800 9520
rect 0 9436 1708 9492
rect 1764 9436 2492 9492
rect 2548 9436 2558 9492
rect 0 9408 800 9436
rect 5126 9380 5136 9436
rect 5192 9380 5240 9436
rect 5296 9380 5344 9436
rect 5400 9380 5410 9436
rect 35846 9380 35856 9436
rect 35912 9380 35960 9436
rect 36016 9380 36064 9436
rect 36120 9380 36130 9436
rect 66566 9380 66576 9436
rect 66632 9380 66680 9436
rect 66736 9380 66784 9436
rect 66840 9380 66850 9436
rect 97286 9380 97296 9436
rect 97352 9380 97400 9436
rect 97456 9380 97504 9436
rect 97560 9380 97570 9436
rect 128006 9380 128016 9436
rect 128072 9380 128120 9436
rect 128176 9380 128224 9436
rect 128280 9380 128290 9436
rect 158726 9380 158736 9436
rect 158792 9380 158840 9436
rect 158896 9380 158944 9436
rect 159000 9380 159010 9436
rect 189446 9380 189456 9436
rect 189512 9380 189560 9436
rect 189616 9380 189664 9436
rect 189720 9380 189730 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 127346 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127630 8652
rect 158066 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158350 8652
rect 188786 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189070 8652
rect 5126 7812 5136 7868
rect 5192 7812 5240 7868
rect 5296 7812 5344 7868
rect 5400 7812 5410 7868
rect 35846 7812 35856 7868
rect 35912 7812 35960 7868
rect 36016 7812 36064 7868
rect 36120 7812 36130 7868
rect 66566 7812 66576 7868
rect 66632 7812 66680 7868
rect 66736 7812 66784 7868
rect 66840 7812 66850 7868
rect 97286 7812 97296 7868
rect 97352 7812 97400 7868
rect 97456 7812 97504 7868
rect 97560 7812 97570 7868
rect 128006 7812 128016 7868
rect 128072 7812 128120 7868
rect 128176 7812 128224 7868
rect 128280 7812 128290 7868
rect 158726 7812 158736 7868
rect 158792 7812 158840 7868
rect 158896 7812 158944 7868
rect 159000 7812 159010 7868
rect 189446 7812 189456 7868
rect 189512 7812 189560 7868
rect 189616 7812 189664 7868
rect 189720 7812 189730 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 127346 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127630 7084
rect 158066 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158350 7084
rect 188786 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189070 7084
rect 5126 6244 5136 6300
rect 5192 6244 5240 6300
rect 5296 6244 5344 6300
rect 5400 6244 5410 6300
rect 35846 6244 35856 6300
rect 35912 6244 35960 6300
rect 36016 6244 36064 6300
rect 36120 6244 36130 6300
rect 66566 6244 66576 6300
rect 66632 6244 66680 6300
rect 66736 6244 66784 6300
rect 66840 6244 66850 6300
rect 97286 6244 97296 6300
rect 97352 6244 97400 6300
rect 97456 6244 97504 6300
rect 97560 6244 97570 6300
rect 128006 6244 128016 6300
rect 128072 6244 128120 6300
rect 128176 6244 128224 6300
rect 128280 6244 128290 6300
rect 158726 6244 158736 6300
rect 158792 6244 158840 6300
rect 158896 6244 158944 6300
rect 159000 6244 159010 6300
rect 189446 6244 189456 6300
rect 189512 6244 189560 6300
rect 189616 6244 189664 6300
rect 189720 6244 189730 6300
rect 0 5684 800 5712
rect 0 5628 1708 5684
rect 1764 5628 1774 5684
rect 0 5600 800 5628
rect 205332 5600 206132 5712
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 127346 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127630 5516
rect 158066 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158350 5516
rect 188786 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189070 5516
rect 5126 4676 5136 4732
rect 5192 4676 5240 4732
rect 5296 4676 5344 4732
rect 5400 4676 5410 4732
rect 35846 4676 35856 4732
rect 35912 4676 35960 4732
rect 36016 4676 36064 4732
rect 36120 4676 36130 4732
rect 66566 4676 66576 4732
rect 66632 4676 66680 4732
rect 66736 4676 66784 4732
rect 66840 4676 66850 4732
rect 97286 4676 97296 4732
rect 97352 4676 97400 4732
rect 97456 4676 97504 4732
rect 97560 4676 97570 4732
rect 128006 4676 128016 4732
rect 128072 4676 128120 4732
rect 128176 4676 128224 4732
rect 128280 4676 128290 4732
rect 158726 4676 158736 4732
rect 158792 4676 158840 4732
rect 158896 4676 158944 4732
rect 159000 4676 159010 4732
rect 189446 4676 189456 4732
rect 189512 4676 189560 4732
rect 189616 4676 189664 4732
rect 189720 4676 189730 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 127346 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127630 3948
rect 158066 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158350 3948
rect 188786 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189070 3948
rect 5126 3108 5136 3164
rect 5192 3108 5240 3164
rect 5296 3108 5344 3164
rect 5400 3108 5410 3164
rect 35846 3108 35856 3164
rect 35912 3108 35960 3164
rect 36016 3108 36064 3164
rect 36120 3108 36130 3164
rect 66566 3108 66576 3164
rect 66632 3108 66680 3164
rect 66736 3108 66784 3164
rect 66840 3108 66850 3164
rect 97286 3108 97296 3164
rect 97352 3108 97400 3164
rect 97456 3108 97504 3164
rect 97560 3108 97570 3164
rect 128006 3108 128016 3164
rect 128072 3108 128120 3164
rect 128176 3108 128224 3164
rect 128280 3108 128290 3164
rect 158726 3108 158736 3164
rect 158792 3108 158840 3164
rect 158896 3108 158944 3164
rect 159000 3108 159010 3164
rect 189446 3108 189456 3164
rect 189512 3108 189560 3164
rect 189616 3108 189664 3164
rect 189720 3108 189730 3164
rect 0 1876 800 1904
rect 0 1820 1708 1876
rect 1764 1820 1774 1876
rect 0 1792 800 1820
<< via3 >>
rect 5136 156772 5192 156828
rect 5240 156772 5296 156828
rect 5344 156772 5400 156828
rect 35856 156772 35912 156828
rect 35960 156772 36016 156828
rect 36064 156772 36120 156828
rect 66576 156772 66632 156828
rect 66680 156772 66736 156828
rect 66784 156772 66840 156828
rect 97296 156772 97352 156828
rect 97400 156772 97456 156828
rect 97504 156772 97560 156828
rect 128016 156772 128072 156828
rect 128120 156772 128176 156828
rect 128224 156772 128280 156828
rect 158736 156772 158792 156828
rect 158840 156772 158896 156828
rect 158944 156772 159000 156828
rect 189456 156772 189512 156828
rect 189560 156772 189616 156828
rect 189664 156772 189720 156828
rect 4476 155988 4532 156044
rect 4580 155988 4636 156044
rect 4684 155988 4740 156044
rect 35196 155988 35252 156044
rect 35300 155988 35356 156044
rect 35404 155988 35460 156044
rect 65916 155988 65972 156044
rect 66020 155988 66076 156044
rect 66124 155988 66180 156044
rect 96636 155988 96692 156044
rect 96740 155988 96796 156044
rect 96844 155988 96900 156044
rect 127356 155988 127412 156044
rect 127460 155988 127516 156044
rect 127564 155988 127620 156044
rect 158076 155988 158132 156044
rect 158180 155988 158236 156044
rect 158284 155988 158340 156044
rect 188796 155988 188852 156044
rect 188900 155988 188956 156044
rect 189004 155988 189060 156044
rect 5136 155204 5192 155260
rect 5240 155204 5296 155260
rect 5344 155204 5400 155260
rect 35856 155204 35912 155260
rect 35960 155204 36016 155260
rect 36064 155204 36120 155260
rect 66576 155204 66632 155260
rect 66680 155204 66736 155260
rect 66784 155204 66840 155260
rect 97296 155204 97352 155260
rect 97400 155204 97456 155260
rect 97504 155204 97560 155260
rect 128016 155204 128072 155260
rect 128120 155204 128176 155260
rect 128224 155204 128280 155260
rect 158736 155204 158792 155260
rect 158840 155204 158896 155260
rect 158944 155204 159000 155260
rect 189456 155204 189512 155260
rect 189560 155204 189616 155260
rect 189664 155204 189720 155260
rect 4476 154420 4532 154476
rect 4580 154420 4636 154476
rect 4684 154420 4740 154476
rect 35196 154420 35252 154476
rect 35300 154420 35356 154476
rect 35404 154420 35460 154476
rect 65916 154420 65972 154476
rect 66020 154420 66076 154476
rect 66124 154420 66180 154476
rect 96636 154420 96692 154476
rect 96740 154420 96796 154476
rect 96844 154420 96900 154476
rect 127356 154420 127412 154476
rect 127460 154420 127516 154476
rect 127564 154420 127620 154476
rect 158076 154420 158132 154476
rect 158180 154420 158236 154476
rect 158284 154420 158340 154476
rect 188796 154420 188852 154476
rect 188900 154420 188956 154476
rect 189004 154420 189060 154476
rect 5136 153636 5192 153692
rect 5240 153636 5296 153692
rect 5344 153636 5400 153692
rect 35856 153636 35912 153692
rect 35960 153636 36016 153692
rect 36064 153636 36120 153692
rect 66576 153636 66632 153692
rect 66680 153636 66736 153692
rect 66784 153636 66840 153692
rect 97296 153636 97352 153692
rect 97400 153636 97456 153692
rect 97504 153636 97560 153692
rect 128016 153636 128072 153692
rect 128120 153636 128176 153692
rect 128224 153636 128280 153692
rect 158736 153636 158792 153692
rect 158840 153636 158896 153692
rect 158944 153636 159000 153692
rect 189456 153636 189512 153692
rect 189560 153636 189616 153692
rect 189664 153636 189720 153692
rect 4476 152852 4532 152908
rect 4580 152852 4636 152908
rect 4684 152852 4740 152908
rect 35196 152852 35252 152908
rect 35300 152852 35356 152908
rect 35404 152852 35460 152908
rect 65916 152852 65972 152908
rect 66020 152852 66076 152908
rect 66124 152852 66180 152908
rect 96636 152852 96692 152908
rect 96740 152852 96796 152908
rect 96844 152852 96900 152908
rect 127356 152852 127412 152908
rect 127460 152852 127516 152908
rect 127564 152852 127620 152908
rect 158076 152852 158132 152908
rect 158180 152852 158236 152908
rect 158284 152852 158340 152908
rect 188796 152852 188852 152908
rect 188900 152852 188956 152908
rect 189004 152852 189060 152908
rect 5136 152068 5192 152124
rect 5240 152068 5296 152124
rect 5344 152068 5400 152124
rect 35856 152068 35912 152124
rect 35960 152068 36016 152124
rect 36064 152068 36120 152124
rect 66576 152068 66632 152124
rect 66680 152068 66736 152124
rect 66784 152068 66840 152124
rect 97296 152068 97352 152124
rect 97400 152068 97456 152124
rect 97504 152068 97560 152124
rect 128016 152068 128072 152124
rect 128120 152068 128176 152124
rect 128224 152068 128280 152124
rect 158736 152068 158792 152124
rect 158840 152068 158896 152124
rect 158944 152068 159000 152124
rect 189456 152068 189512 152124
rect 189560 152068 189616 152124
rect 189664 152068 189720 152124
rect 4476 151284 4532 151340
rect 4580 151284 4636 151340
rect 4684 151284 4740 151340
rect 35196 151284 35252 151340
rect 35300 151284 35356 151340
rect 35404 151284 35460 151340
rect 65916 151284 65972 151340
rect 66020 151284 66076 151340
rect 66124 151284 66180 151340
rect 96636 151284 96692 151340
rect 96740 151284 96796 151340
rect 96844 151284 96900 151340
rect 127356 151284 127412 151340
rect 127460 151284 127516 151340
rect 127564 151284 127620 151340
rect 158076 151284 158132 151340
rect 158180 151284 158236 151340
rect 158284 151284 158340 151340
rect 188796 151284 188852 151340
rect 188900 151284 188956 151340
rect 189004 151284 189060 151340
rect 5136 150500 5192 150556
rect 5240 150500 5296 150556
rect 5344 150500 5400 150556
rect 35856 150500 35912 150556
rect 35960 150500 36016 150556
rect 36064 150500 36120 150556
rect 66576 150500 66632 150556
rect 66680 150500 66736 150556
rect 66784 150500 66840 150556
rect 97296 150500 97352 150556
rect 97400 150500 97456 150556
rect 97504 150500 97560 150556
rect 128016 150500 128072 150556
rect 128120 150500 128176 150556
rect 128224 150500 128280 150556
rect 158736 150500 158792 150556
rect 158840 150500 158896 150556
rect 158944 150500 159000 150556
rect 189456 150500 189512 150556
rect 189560 150500 189616 150556
rect 189664 150500 189720 150556
rect 4476 149716 4532 149772
rect 4580 149716 4636 149772
rect 4684 149716 4740 149772
rect 35196 149716 35252 149772
rect 35300 149716 35356 149772
rect 35404 149716 35460 149772
rect 65916 149716 65972 149772
rect 66020 149716 66076 149772
rect 66124 149716 66180 149772
rect 96636 149716 96692 149772
rect 96740 149716 96796 149772
rect 96844 149716 96900 149772
rect 127356 149716 127412 149772
rect 127460 149716 127516 149772
rect 127564 149716 127620 149772
rect 158076 149716 158132 149772
rect 158180 149716 158236 149772
rect 158284 149716 158340 149772
rect 188796 149716 188852 149772
rect 188900 149716 188956 149772
rect 189004 149716 189060 149772
rect 5136 148932 5192 148988
rect 5240 148932 5296 148988
rect 5344 148932 5400 148988
rect 35856 148932 35912 148988
rect 35960 148932 36016 148988
rect 36064 148932 36120 148988
rect 66576 148932 66632 148988
rect 66680 148932 66736 148988
rect 66784 148932 66840 148988
rect 97296 148932 97352 148988
rect 97400 148932 97456 148988
rect 97504 148932 97560 148988
rect 128016 148932 128072 148988
rect 128120 148932 128176 148988
rect 128224 148932 128280 148988
rect 158736 148932 158792 148988
rect 158840 148932 158896 148988
rect 158944 148932 159000 148988
rect 189456 148932 189512 148988
rect 189560 148932 189616 148988
rect 189664 148932 189720 148988
rect 4476 148148 4532 148204
rect 4580 148148 4636 148204
rect 4684 148148 4740 148204
rect 35196 148148 35252 148204
rect 35300 148148 35356 148204
rect 35404 148148 35460 148204
rect 65916 148148 65972 148204
rect 66020 148148 66076 148204
rect 66124 148148 66180 148204
rect 96636 148148 96692 148204
rect 96740 148148 96796 148204
rect 96844 148148 96900 148204
rect 127356 148148 127412 148204
rect 127460 148148 127516 148204
rect 127564 148148 127620 148204
rect 158076 148148 158132 148204
rect 158180 148148 158236 148204
rect 158284 148148 158340 148204
rect 188796 148148 188852 148204
rect 188900 148148 188956 148204
rect 189004 148148 189060 148204
rect 5136 147364 5192 147420
rect 5240 147364 5296 147420
rect 5344 147364 5400 147420
rect 35856 147364 35912 147420
rect 35960 147364 36016 147420
rect 36064 147364 36120 147420
rect 66576 147364 66632 147420
rect 66680 147364 66736 147420
rect 66784 147364 66840 147420
rect 97296 147364 97352 147420
rect 97400 147364 97456 147420
rect 97504 147364 97560 147420
rect 128016 147364 128072 147420
rect 128120 147364 128176 147420
rect 128224 147364 128280 147420
rect 158736 147364 158792 147420
rect 158840 147364 158896 147420
rect 158944 147364 159000 147420
rect 189456 147364 189512 147420
rect 189560 147364 189616 147420
rect 189664 147364 189720 147420
rect 4476 146580 4532 146636
rect 4580 146580 4636 146636
rect 4684 146580 4740 146636
rect 35196 146580 35252 146636
rect 35300 146580 35356 146636
rect 35404 146580 35460 146636
rect 65916 146580 65972 146636
rect 66020 146580 66076 146636
rect 66124 146580 66180 146636
rect 96636 146580 96692 146636
rect 96740 146580 96796 146636
rect 96844 146580 96900 146636
rect 127356 146580 127412 146636
rect 127460 146580 127516 146636
rect 127564 146580 127620 146636
rect 158076 146580 158132 146636
rect 158180 146580 158236 146636
rect 158284 146580 158340 146636
rect 188796 146580 188852 146636
rect 188900 146580 188956 146636
rect 189004 146580 189060 146636
rect 5136 145796 5192 145852
rect 5240 145796 5296 145852
rect 5344 145796 5400 145852
rect 35856 145796 35912 145852
rect 35960 145796 36016 145852
rect 36064 145796 36120 145852
rect 66576 145796 66632 145852
rect 66680 145796 66736 145852
rect 66784 145796 66840 145852
rect 97296 145796 97352 145852
rect 97400 145796 97456 145852
rect 97504 145796 97560 145852
rect 128016 145796 128072 145852
rect 128120 145796 128176 145852
rect 128224 145796 128280 145852
rect 158736 145796 158792 145852
rect 158840 145796 158896 145852
rect 158944 145796 159000 145852
rect 189456 145796 189512 145852
rect 189560 145796 189616 145852
rect 189664 145796 189720 145852
rect 4476 145012 4532 145068
rect 4580 145012 4636 145068
rect 4684 145012 4740 145068
rect 35196 145012 35252 145068
rect 35300 145012 35356 145068
rect 35404 145012 35460 145068
rect 65916 145012 65972 145068
rect 66020 145012 66076 145068
rect 66124 145012 66180 145068
rect 96636 145012 96692 145068
rect 96740 145012 96796 145068
rect 96844 145012 96900 145068
rect 127356 145012 127412 145068
rect 127460 145012 127516 145068
rect 127564 145012 127620 145068
rect 158076 145012 158132 145068
rect 158180 145012 158236 145068
rect 158284 145012 158340 145068
rect 188796 145012 188852 145068
rect 188900 145012 188956 145068
rect 189004 145012 189060 145068
rect 5136 144228 5192 144284
rect 5240 144228 5296 144284
rect 5344 144228 5400 144284
rect 189456 144228 189512 144284
rect 189560 144228 189616 144284
rect 189664 144228 189720 144284
rect 4476 143444 4532 143500
rect 4580 143444 4636 143500
rect 4684 143444 4740 143500
rect 188796 143444 188852 143500
rect 188900 143444 188956 143500
rect 189004 143444 189060 143500
rect 5136 142660 5192 142716
rect 5240 142660 5296 142716
rect 5344 142660 5400 142716
rect 189456 142660 189512 142716
rect 189560 142660 189616 142716
rect 189664 142660 189720 142716
rect 4476 141876 4532 141932
rect 4580 141876 4636 141932
rect 4684 141876 4740 141932
rect 188796 141876 188852 141932
rect 188900 141876 188956 141932
rect 189004 141876 189060 141932
rect 5136 141092 5192 141148
rect 5240 141092 5296 141148
rect 5344 141092 5400 141148
rect 189456 141092 189512 141148
rect 189560 141092 189616 141148
rect 189664 141092 189720 141148
rect 4476 140308 4532 140364
rect 4580 140308 4636 140364
rect 4684 140308 4740 140364
rect 188796 140308 188852 140364
rect 188900 140308 188956 140364
rect 189004 140308 189060 140364
rect 5136 139524 5192 139580
rect 5240 139524 5296 139580
rect 5344 139524 5400 139580
rect 189456 139524 189512 139580
rect 189560 139524 189616 139580
rect 189664 139524 189720 139580
rect 4476 138740 4532 138796
rect 4580 138740 4636 138796
rect 4684 138740 4740 138796
rect 188796 138740 188852 138796
rect 188900 138740 188956 138796
rect 189004 138740 189060 138796
rect 5136 137956 5192 138012
rect 5240 137956 5296 138012
rect 5344 137956 5400 138012
rect 189456 137956 189512 138012
rect 189560 137956 189616 138012
rect 189664 137956 189720 138012
rect 4476 137172 4532 137228
rect 4580 137172 4636 137228
rect 4684 137172 4740 137228
rect 188796 137172 188852 137228
rect 188900 137172 188956 137228
rect 189004 137172 189060 137228
rect 5136 136388 5192 136444
rect 5240 136388 5296 136444
rect 5344 136388 5400 136444
rect 189456 136388 189512 136444
rect 189560 136388 189616 136444
rect 189664 136388 189720 136444
rect 4476 135604 4532 135660
rect 4580 135604 4636 135660
rect 4684 135604 4740 135660
rect 188796 135604 188852 135660
rect 188900 135604 188956 135660
rect 189004 135604 189060 135660
rect 5136 134820 5192 134876
rect 5240 134820 5296 134876
rect 5344 134820 5400 134876
rect 189456 134820 189512 134876
rect 189560 134820 189616 134876
rect 189664 134820 189720 134876
rect 4476 134036 4532 134092
rect 4580 134036 4636 134092
rect 4684 134036 4740 134092
rect 188796 134036 188852 134092
rect 188900 134036 188956 134092
rect 189004 134036 189060 134092
rect 5136 133252 5192 133308
rect 5240 133252 5296 133308
rect 5344 133252 5400 133308
rect 189456 133252 189512 133308
rect 189560 133252 189616 133308
rect 189664 133252 189720 133308
rect 4476 132468 4532 132524
rect 4580 132468 4636 132524
rect 4684 132468 4740 132524
rect 188796 132468 188852 132524
rect 188900 132468 188956 132524
rect 189004 132468 189060 132524
rect 5136 131684 5192 131740
rect 5240 131684 5296 131740
rect 5344 131684 5400 131740
rect 189456 131684 189512 131740
rect 189560 131684 189616 131740
rect 189664 131684 189720 131740
rect 4476 130900 4532 130956
rect 4580 130900 4636 130956
rect 4684 130900 4740 130956
rect 188796 130900 188852 130956
rect 188900 130900 188956 130956
rect 189004 130900 189060 130956
rect 5136 130116 5192 130172
rect 5240 130116 5296 130172
rect 5344 130116 5400 130172
rect 189456 130116 189512 130172
rect 189560 130116 189616 130172
rect 189664 130116 189720 130172
rect 4476 129332 4532 129388
rect 4580 129332 4636 129388
rect 4684 129332 4740 129388
rect 188796 129332 188852 129388
rect 188900 129332 188956 129388
rect 189004 129332 189060 129388
rect 5136 128548 5192 128604
rect 5240 128548 5296 128604
rect 5344 128548 5400 128604
rect 189456 128548 189512 128604
rect 189560 128548 189616 128604
rect 189664 128548 189720 128604
rect 4476 127764 4532 127820
rect 4580 127764 4636 127820
rect 4684 127764 4740 127820
rect 188796 127764 188852 127820
rect 188900 127764 188956 127820
rect 189004 127764 189060 127820
rect 5136 126980 5192 127036
rect 5240 126980 5296 127036
rect 5344 126980 5400 127036
rect 189456 126980 189512 127036
rect 189560 126980 189616 127036
rect 189664 126980 189720 127036
rect 4476 126196 4532 126252
rect 4580 126196 4636 126252
rect 4684 126196 4740 126252
rect 188796 126196 188852 126252
rect 188900 126196 188956 126252
rect 189004 126196 189060 126252
rect 5136 125412 5192 125468
rect 5240 125412 5296 125468
rect 5344 125412 5400 125468
rect 189456 125412 189512 125468
rect 189560 125412 189616 125468
rect 189664 125412 189720 125468
rect 4476 124628 4532 124684
rect 4580 124628 4636 124684
rect 4684 124628 4740 124684
rect 188796 124628 188852 124684
rect 188900 124628 188956 124684
rect 189004 124628 189060 124684
rect 5136 123844 5192 123900
rect 5240 123844 5296 123900
rect 5344 123844 5400 123900
rect 189456 123844 189512 123900
rect 189560 123844 189616 123900
rect 189664 123844 189720 123900
rect 4476 123060 4532 123116
rect 4580 123060 4636 123116
rect 4684 123060 4740 123116
rect 188796 123060 188852 123116
rect 188900 123060 188956 123116
rect 189004 123060 189060 123116
rect 5136 122276 5192 122332
rect 5240 122276 5296 122332
rect 5344 122276 5400 122332
rect 189456 122276 189512 122332
rect 189560 122276 189616 122332
rect 189664 122276 189720 122332
rect 4476 121492 4532 121548
rect 4580 121492 4636 121548
rect 4684 121492 4740 121548
rect 188796 121492 188852 121548
rect 188900 121492 188956 121548
rect 189004 121492 189060 121548
rect 5136 120708 5192 120764
rect 5240 120708 5296 120764
rect 5344 120708 5400 120764
rect 189456 120708 189512 120764
rect 189560 120708 189616 120764
rect 189664 120708 189720 120764
rect 4476 119924 4532 119980
rect 4580 119924 4636 119980
rect 4684 119924 4740 119980
rect 188796 119924 188852 119980
rect 188900 119924 188956 119980
rect 189004 119924 189060 119980
rect 5136 119140 5192 119196
rect 5240 119140 5296 119196
rect 5344 119140 5400 119196
rect 189456 119140 189512 119196
rect 189560 119140 189616 119196
rect 189664 119140 189720 119196
rect 4476 118356 4532 118412
rect 4580 118356 4636 118412
rect 4684 118356 4740 118412
rect 188796 118356 188852 118412
rect 188900 118356 188956 118412
rect 189004 118356 189060 118412
rect 5136 117572 5192 117628
rect 5240 117572 5296 117628
rect 5344 117572 5400 117628
rect 189456 117572 189512 117628
rect 189560 117572 189616 117628
rect 189664 117572 189720 117628
rect 4476 116788 4532 116844
rect 4580 116788 4636 116844
rect 4684 116788 4740 116844
rect 188796 116788 188852 116844
rect 188900 116788 188956 116844
rect 189004 116788 189060 116844
rect 5136 116004 5192 116060
rect 5240 116004 5296 116060
rect 5344 116004 5400 116060
rect 189456 116004 189512 116060
rect 189560 116004 189616 116060
rect 189664 116004 189720 116060
rect 4476 115220 4532 115276
rect 4580 115220 4636 115276
rect 4684 115220 4740 115276
rect 188796 115220 188852 115276
rect 188900 115220 188956 115276
rect 189004 115220 189060 115276
rect 5136 114436 5192 114492
rect 5240 114436 5296 114492
rect 5344 114436 5400 114492
rect 189456 114436 189512 114492
rect 189560 114436 189616 114492
rect 189664 114436 189720 114492
rect 4476 113652 4532 113708
rect 4580 113652 4636 113708
rect 4684 113652 4740 113708
rect 188796 113652 188852 113708
rect 188900 113652 188956 113708
rect 189004 113652 189060 113708
rect 5136 112868 5192 112924
rect 5240 112868 5296 112924
rect 5344 112868 5400 112924
rect 189456 112868 189512 112924
rect 189560 112868 189616 112924
rect 189664 112868 189720 112924
rect 4476 112084 4532 112140
rect 4580 112084 4636 112140
rect 4684 112084 4740 112140
rect 188796 112084 188852 112140
rect 188900 112084 188956 112140
rect 189004 112084 189060 112140
rect 5136 111300 5192 111356
rect 5240 111300 5296 111356
rect 5344 111300 5400 111356
rect 189456 111300 189512 111356
rect 189560 111300 189616 111356
rect 189664 111300 189720 111356
rect 4476 110516 4532 110572
rect 4580 110516 4636 110572
rect 4684 110516 4740 110572
rect 188796 110516 188852 110572
rect 188900 110516 188956 110572
rect 189004 110516 189060 110572
rect 5136 109732 5192 109788
rect 5240 109732 5296 109788
rect 5344 109732 5400 109788
rect 189456 109732 189512 109788
rect 189560 109732 189616 109788
rect 189664 109732 189720 109788
rect 4476 108948 4532 109004
rect 4580 108948 4636 109004
rect 4684 108948 4740 109004
rect 188796 108948 188852 109004
rect 188900 108948 188956 109004
rect 189004 108948 189060 109004
rect 5136 108164 5192 108220
rect 5240 108164 5296 108220
rect 5344 108164 5400 108220
rect 189456 108164 189512 108220
rect 189560 108164 189616 108220
rect 189664 108164 189720 108220
rect 4476 107380 4532 107436
rect 4580 107380 4636 107436
rect 4684 107380 4740 107436
rect 188796 107380 188852 107436
rect 188900 107380 188956 107436
rect 189004 107380 189060 107436
rect 5136 106596 5192 106652
rect 5240 106596 5296 106652
rect 5344 106596 5400 106652
rect 189456 106596 189512 106652
rect 189560 106596 189616 106652
rect 189664 106596 189720 106652
rect 4476 105812 4532 105868
rect 4580 105812 4636 105868
rect 4684 105812 4740 105868
rect 188796 105812 188852 105868
rect 188900 105812 188956 105868
rect 189004 105812 189060 105868
rect 5136 105028 5192 105084
rect 5240 105028 5296 105084
rect 5344 105028 5400 105084
rect 189456 105028 189512 105084
rect 189560 105028 189616 105084
rect 189664 105028 189720 105084
rect 4476 104244 4532 104300
rect 4580 104244 4636 104300
rect 4684 104244 4740 104300
rect 188796 104244 188852 104300
rect 188900 104244 188956 104300
rect 189004 104244 189060 104300
rect 5136 103460 5192 103516
rect 5240 103460 5296 103516
rect 5344 103460 5400 103516
rect 189456 103460 189512 103516
rect 189560 103460 189616 103516
rect 189664 103460 189720 103516
rect 4476 102676 4532 102732
rect 4580 102676 4636 102732
rect 4684 102676 4740 102732
rect 188796 102676 188852 102732
rect 188900 102676 188956 102732
rect 189004 102676 189060 102732
rect 5136 101892 5192 101948
rect 5240 101892 5296 101948
rect 5344 101892 5400 101948
rect 189456 101892 189512 101948
rect 189560 101892 189616 101948
rect 189664 101892 189720 101948
rect 4476 101108 4532 101164
rect 4580 101108 4636 101164
rect 4684 101108 4740 101164
rect 188796 101108 188852 101164
rect 188900 101108 188956 101164
rect 189004 101108 189060 101164
rect 5136 100324 5192 100380
rect 5240 100324 5296 100380
rect 5344 100324 5400 100380
rect 189456 100324 189512 100380
rect 189560 100324 189616 100380
rect 189664 100324 189720 100380
rect 4476 99540 4532 99596
rect 4580 99540 4636 99596
rect 4684 99540 4740 99596
rect 188796 99540 188852 99596
rect 188900 99540 188956 99596
rect 189004 99540 189060 99596
rect 5136 98756 5192 98812
rect 5240 98756 5296 98812
rect 5344 98756 5400 98812
rect 189456 98756 189512 98812
rect 189560 98756 189616 98812
rect 189664 98756 189720 98812
rect 4476 97972 4532 98028
rect 4580 97972 4636 98028
rect 4684 97972 4740 98028
rect 188796 97972 188852 98028
rect 188900 97972 188956 98028
rect 189004 97972 189060 98028
rect 5136 97188 5192 97244
rect 5240 97188 5296 97244
rect 5344 97188 5400 97244
rect 189456 97188 189512 97244
rect 189560 97188 189616 97244
rect 189664 97188 189720 97244
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 188796 96404 188852 96460
rect 188900 96404 188956 96460
rect 189004 96404 189060 96460
rect 5136 95620 5192 95676
rect 5240 95620 5296 95676
rect 5344 95620 5400 95676
rect 189456 95620 189512 95676
rect 189560 95620 189616 95676
rect 189664 95620 189720 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 188796 94836 188852 94892
rect 188900 94836 188956 94892
rect 189004 94836 189060 94892
rect 5136 94052 5192 94108
rect 5240 94052 5296 94108
rect 5344 94052 5400 94108
rect 189456 94052 189512 94108
rect 189560 94052 189616 94108
rect 189664 94052 189720 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 188796 93268 188852 93324
rect 188900 93268 188956 93324
rect 189004 93268 189060 93324
rect 5136 92484 5192 92540
rect 5240 92484 5296 92540
rect 5344 92484 5400 92540
rect 189456 92484 189512 92540
rect 189560 92484 189616 92540
rect 189664 92484 189720 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 188796 91700 188852 91756
rect 188900 91700 188956 91756
rect 189004 91700 189060 91756
rect 5136 90916 5192 90972
rect 5240 90916 5296 90972
rect 5344 90916 5400 90972
rect 189456 90916 189512 90972
rect 189560 90916 189616 90972
rect 189664 90916 189720 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 188796 90132 188852 90188
rect 188900 90132 188956 90188
rect 189004 90132 189060 90188
rect 5136 89348 5192 89404
rect 5240 89348 5296 89404
rect 5344 89348 5400 89404
rect 189456 89348 189512 89404
rect 189560 89348 189616 89404
rect 189664 89348 189720 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 188796 88564 188852 88620
rect 188900 88564 188956 88620
rect 189004 88564 189060 88620
rect 5136 87780 5192 87836
rect 5240 87780 5296 87836
rect 5344 87780 5400 87836
rect 189456 87780 189512 87836
rect 189560 87780 189616 87836
rect 189664 87780 189720 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 188796 86996 188852 87052
rect 188900 86996 188956 87052
rect 189004 86996 189060 87052
rect 5136 86212 5192 86268
rect 5240 86212 5296 86268
rect 5344 86212 5400 86268
rect 189456 86212 189512 86268
rect 189560 86212 189616 86268
rect 189664 86212 189720 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 188796 85428 188852 85484
rect 188900 85428 188956 85484
rect 189004 85428 189060 85484
rect 5136 84644 5192 84700
rect 5240 84644 5296 84700
rect 5344 84644 5400 84700
rect 189456 84644 189512 84700
rect 189560 84644 189616 84700
rect 189664 84644 189720 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 188796 83860 188852 83916
rect 188900 83860 188956 83916
rect 189004 83860 189060 83916
rect 5136 83076 5192 83132
rect 5240 83076 5296 83132
rect 5344 83076 5400 83132
rect 189456 83076 189512 83132
rect 189560 83076 189616 83132
rect 189664 83076 189720 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 188796 82292 188852 82348
rect 188900 82292 188956 82348
rect 189004 82292 189060 82348
rect 5136 81508 5192 81564
rect 5240 81508 5296 81564
rect 5344 81508 5400 81564
rect 189456 81508 189512 81564
rect 189560 81508 189616 81564
rect 189664 81508 189720 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 188796 80724 188852 80780
rect 188900 80724 188956 80780
rect 189004 80724 189060 80780
rect 5136 79940 5192 79996
rect 5240 79940 5296 79996
rect 5344 79940 5400 79996
rect 189456 79940 189512 79996
rect 189560 79940 189616 79996
rect 189664 79940 189720 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 188796 79156 188852 79212
rect 188900 79156 188956 79212
rect 189004 79156 189060 79212
rect 5136 78372 5192 78428
rect 5240 78372 5296 78428
rect 5344 78372 5400 78428
rect 189456 78372 189512 78428
rect 189560 78372 189616 78428
rect 189664 78372 189720 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 188796 77588 188852 77644
rect 188900 77588 188956 77644
rect 189004 77588 189060 77644
rect 5136 76804 5192 76860
rect 5240 76804 5296 76860
rect 5344 76804 5400 76860
rect 189456 76804 189512 76860
rect 189560 76804 189616 76860
rect 189664 76804 189720 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 188796 76020 188852 76076
rect 188900 76020 188956 76076
rect 189004 76020 189060 76076
rect 5136 75236 5192 75292
rect 5240 75236 5296 75292
rect 5344 75236 5400 75292
rect 189456 75236 189512 75292
rect 189560 75236 189616 75292
rect 189664 75236 189720 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 188796 74452 188852 74508
rect 188900 74452 188956 74508
rect 189004 74452 189060 74508
rect 5136 73668 5192 73724
rect 5240 73668 5296 73724
rect 5344 73668 5400 73724
rect 189456 73668 189512 73724
rect 189560 73668 189616 73724
rect 189664 73668 189720 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 188796 72884 188852 72940
rect 188900 72884 188956 72940
rect 189004 72884 189060 72940
rect 5136 72100 5192 72156
rect 5240 72100 5296 72156
rect 5344 72100 5400 72156
rect 189456 72100 189512 72156
rect 189560 72100 189616 72156
rect 189664 72100 189720 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 188796 71316 188852 71372
rect 188900 71316 188956 71372
rect 189004 71316 189060 71372
rect 5136 70532 5192 70588
rect 5240 70532 5296 70588
rect 5344 70532 5400 70588
rect 189456 70532 189512 70588
rect 189560 70532 189616 70588
rect 189664 70532 189720 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 188796 69748 188852 69804
rect 188900 69748 188956 69804
rect 189004 69748 189060 69804
rect 5136 68964 5192 69020
rect 5240 68964 5296 69020
rect 5344 68964 5400 69020
rect 189456 68964 189512 69020
rect 189560 68964 189616 69020
rect 189664 68964 189720 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 188796 68180 188852 68236
rect 188900 68180 188956 68236
rect 189004 68180 189060 68236
rect 5136 67396 5192 67452
rect 5240 67396 5296 67452
rect 5344 67396 5400 67452
rect 189456 67396 189512 67452
rect 189560 67396 189616 67452
rect 189664 67396 189720 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 188796 66612 188852 66668
rect 188900 66612 188956 66668
rect 189004 66612 189060 66668
rect 5136 65828 5192 65884
rect 5240 65828 5296 65884
rect 5344 65828 5400 65884
rect 189456 65828 189512 65884
rect 189560 65828 189616 65884
rect 189664 65828 189720 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 188796 65044 188852 65100
rect 188900 65044 188956 65100
rect 189004 65044 189060 65100
rect 5136 64260 5192 64316
rect 5240 64260 5296 64316
rect 5344 64260 5400 64316
rect 189456 64260 189512 64316
rect 189560 64260 189616 64316
rect 189664 64260 189720 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 188796 63476 188852 63532
rect 188900 63476 188956 63532
rect 189004 63476 189060 63532
rect 5136 62692 5192 62748
rect 5240 62692 5296 62748
rect 5344 62692 5400 62748
rect 189456 62692 189512 62748
rect 189560 62692 189616 62748
rect 189664 62692 189720 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 188796 61908 188852 61964
rect 188900 61908 188956 61964
rect 189004 61908 189060 61964
rect 5136 61124 5192 61180
rect 5240 61124 5296 61180
rect 5344 61124 5400 61180
rect 189456 61124 189512 61180
rect 189560 61124 189616 61180
rect 189664 61124 189720 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 188796 60340 188852 60396
rect 188900 60340 188956 60396
rect 189004 60340 189060 60396
rect 5136 59556 5192 59612
rect 5240 59556 5296 59612
rect 5344 59556 5400 59612
rect 189456 59556 189512 59612
rect 189560 59556 189616 59612
rect 189664 59556 189720 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 188796 58772 188852 58828
rect 188900 58772 188956 58828
rect 189004 58772 189060 58828
rect 5136 57988 5192 58044
rect 5240 57988 5296 58044
rect 5344 57988 5400 58044
rect 189456 57988 189512 58044
rect 189560 57988 189616 58044
rect 189664 57988 189720 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 188796 57204 188852 57260
rect 188900 57204 188956 57260
rect 189004 57204 189060 57260
rect 5136 56420 5192 56476
rect 5240 56420 5296 56476
rect 5344 56420 5400 56476
rect 189456 56420 189512 56476
rect 189560 56420 189616 56476
rect 189664 56420 189720 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 188796 55636 188852 55692
rect 188900 55636 188956 55692
rect 189004 55636 189060 55692
rect 5136 54852 5192 54908
rect 5240 54852 5296 54908
rect 5344 54852 5400 54908
rect 189456 54852 189512 54908
rect 189560 54852 189616 54908
rect 189664 54852 189720 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 188796 54068 188852 54124
rect 188900 54068 188956 54124
rect 189004 54068 189060 54124
rect 5136 53284 5192 53340
rect 5240 53284 5296 53340
rect 5344 53284 5400 53340
rect 189456 53284 189512 53340
rect 189560 53284 189616 53340
rect 189664 53284 189720 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 188796 52500 188852 52556
rect 188900 52500 188956 52556
rect 189004 52500 189060 52556
rect 5136 51716 5192 51772
rect 5240 51716 5296 51772
rect 5344 51716 5400 51772
rect 189456 51716 189512 51772
rect 189560 51716 189616 51772
rect 189664 51716 189720 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 188796 50932 188852 50988
rect 188900 50932 188956 50988
rect 189004 50932 189060 50988
rect 5136 50148 5192 50204
rect 5240 50148 5296 50204
rect 5344 50148 5400 50204
rect 189456 50148 189512 50204
rect 189560 50148 189616 50204
rect 189664 50148 189720 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 188796 49364 188852 49420
rect 188900 49364 188956 49420
rect 189004 49364 189060 49420
rect 5136 48580 5192 48636
rect 5240 48580 5296 48636
rect 5344 48580 5400 48636
rect 189456 48580 189512 48636
rect 189560 48580 189616 48636
rect 189664 48580 189720 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 188796 47796 188852 47852
rect 188900 47796 188956 47852
rect 189004 47796 189060 47852
rect 5136 47012 5192 47068
rect 5240 47012 5296 47068
rect 5344 47012 5400 47068
rect 189456 47012 189512 47068
rect 189560 47012 189616 47068
rect 189664 47012 189720 47068
rect 132972 46956 133028 47012
rect 156380 46956 156436 47012
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 188796 46228 188852 46284
rect 188900 46228 188956 46284
rect 189004 46228 189060 46284
rect 132972 45724 133028 45780
rect 156380 45724 156436 45780
rect 5136 45444 5192 45500
rect 5240 45444 5296 45500
rect 5344 45444 5400 45500
rect 189456 45444 189512 45500
rect 189560 45444 189616 45500
rect 189664 45444 189720 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 188796 44660 188852 44716
rect 188900 44660 188956 44716
rect 189004 44660 189060 44716
rect 5136 43876 5192 43932
rect 5240 43876 5296 43932
rect 5344 43876 5400 43932
rect 189456 43876 189512 43932
rect 189560 43876 189616 43932
rect 189664 43876 189720 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 188796 43092 188852 43148
rect 188900 43092 188956 43148
rect 189004 43092 189060 43148
rect 5136 42308 5192 42364
rect 5240 42308 5296 42364
rect 5344 42308 5400 42364
rect 189456 42308 189512 42364
rect 189560 42308 189616 42364
rect 189664 42308 189720 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 188796 41524 188852 41580
rect 188900 41524 188956 41580
rect 189004 41524 189060 41580
rect 5136 40740 5192 40796
rect 5240 40740 5296 40796
rect 5344 40740 5400 40796
rect 189456 40740 189512 40796
rect 189560 40740 189616 40796
rect 189664 40740 189720 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 188796 39956 188852 40012
rect 188900 39956 188956 40012
rect 189004 39956 189060 40012
rect 5136 39172 5192 39228
rect 5240 39172 5296 39228
rect 5344 39172 5400 39228
rect 189456 39172 189512 39228
rect 189560 39172 189616 39228
rect 189664 39172 189720 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 188796 38388 188852 38444
rect 188900 38388 188956 38444
rect 189004 38388 189060 38444
rect 5136 37604 5192 37660
rect 5240 37604 5296 37660
rect 5344 37604 5400 37660
rect 189456 37604 189512 37660
rect 189560 37604 189616 37660
rect 189664 37604 189720 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 188796 36820 188852 36876
rect 188900 36820 188956 36876
rect 189004 36820 189060 36876
rect 5136 36036 5192 36092
rect 5240 36036 5296 36092
rect 5344 36036 5400 36092
rect 189456 36036 189512 36092
rect 189560 36036 189616 36092
rect 189664 36036 189720 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 188796 35252 188852 35308
rect 188900 35252 188956 35308
rect 189004 35252 189060 35308
rect 5136 34468 5192 34524
rect 5240 34468 5296 34524
rect 5344 34468 5400 34524
rect 189456 34468 189512 34524
rect 189560 34468 189616 34524
rect 189664 34468 189720 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 188796 33684 188852 33740
rect 188900 33684 188956 33740
rect 189004 33684 189060 33740
rect 5136 32900 5192 32956
rect 5240 32900 5296 32956
rect 5344 32900 5400 32956
rect 189456 32900 189512 32956
rect 189560 32900 189616 32956
rect 189664 32900 189720 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 188796 32116 188852 32172
rect 188900 32116 188956 32172
rect 189004 32116 189060 32172
rect 82348 31836 82404 31892
rect 5136 31332 5192 31388
rect 5240 31332 5296 31388
rect 5344 31332 5400 31388
rect 189456 31332 189512 31388
rect 189560 31332 189616 31388
rect 189664 31332 189720 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 188796 30548 188852 30604
rect 188900 30548 188956 30604
rect 189004 30548 189060 30604
rect 5136 29764 5192 29820
rect 5240 29764 5296 29820
rect 5344 29764 5400 29820
rect 189456 29764 189512 29820
rect 189560 29764 189616 29820
rect 189664 29764 189720 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 188796 28980 188852 29036
rect 188900 28980 188956 29036
rect 189004 28980 189060 29036
rect 5136 28196 5192 28252
rect 5240 28196 5296 28252
rect 5344 28196 5400 28252
rect 189456 28196 189512 28252
rect 189560 28196 189616 28252
rect 189664 28196 189720 28252
rect 154700 27804 154756 27860
rect 155148 27692 155204 27748
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 188796 27412 188852 27468
rect 188900 27412 188956 27468
rect 189004 27412 189060 27468
rect 5136 26628 5192 26684
rect 5240 26628 5296 26684
rect 5344 26628 5400 26684
rect 189456 26628 189512 26684
rect 189560 26628 189616 26684
rect 189664 26628 189720 26684
rect 140028 26124 140084 26180
rect 154700 26124 154756 26180
rect 125356 26012 125412 26068
rect 154812 26012 154868 26068
rect 155148 26012 155204 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 188796 25844 188852 25900
rect 188900 25844 188956 25900
rect 189004 25844 189060 25900
rect 96572 25452 96628 25508
rect 77196 25340 77252 25396
rect 110908 25340 110964 25396
rect 78652 25228 78708 25284
rect 82012 25228 82068 25284
rect 5136 25060 5192 25116
rect 5240 25060 5296 25116
rect 5344 25060 5400 25116
rect 189456 25060 189512 25116
rect 189560 25060 189616 25116
rect 189664 25060 189720 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 188796 24276 188852 24332
rect 188900 24276 188956 24332
rect 189004 24276 189060 24332
rect 5136 23492 5192 23548
rect 5240 23492 5296 23548
rect 5344 23492 5400 23548
rect 189456 23492 189512 23548
rect 189560 23492 189616 23548
rect 189664 23492 189720 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 188796 22708 188852 22764
rect 188900 22708 188956 22764
rect 189004 22708 189060 22764
rect 5136 21924 5192 21980
rect 5240 21924 5296 21980
rect 5344 21924 5400 21980
rect 189456 21924 189512 21980
rect 189560 21924 189616 21980
rect 189664 21924 189720 21980
rect 44156 21756 44212 21812
rect 54348 21756 54404 21812
rect 68348 21756 68404 21812
rect 75292 21756 75348 21812
rect 55132 21644 55188 21700
rect 44716 21196 44772 21252
rect 78652 21196 78708 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 188796 21140 188852 21196
rect 188900 21140 188956 21196
rect 189004 21140 189060 21196
rect 77196 21084 77252 21140
rect 48300 20412 48356 20468
rect 67788 20412 67844 20468
rect 82460 20412 82516 20468
rect 154252 20412 154308 20468
rect 5136 20356 5192 20412
rect 5240 20356 5296 20412
rect 5344 20356 5400 20412
rect 189456 20356 189512 20412
rect 189560 20356 189616 20412
rect 189664 20356 189720 20412
rect 58716 19852 58772 19908
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 188796 19572 188852 19628
rect 188900 19572 188956 19628
rect 189004 19572 189060 19628
rect 5136 18788 5192 18844
rect 5240 18788 5296 18844
rect 5344 18788 5400 18844
rect 189456 18788 189512 18844
rect 189560 18788 189616 18844
rect 189664 18788 189720 18844
rect 77308 18396 77364 18452
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 188796 18004 188852 18060
rect 188900 18004 188956 18060
rect 189004 18004 189060 18060
rect 5136 17220 5192 17276
rect 5240 17220 5296 17276
rect 5344 17220 5400 17276
rect 35856 17220 35912 17276
rect 35960 17220 36016 17276
rect 36064 17220 36120 17276
rect 66576 17220 66632 17276
rect 66680 17220 66736 17276
rect 66784 17220 66840 17276
rect 97296 17220 97352 17276
rect 97400 17220 97456 17276
rect 97504 17220 97560 17276
rect 128016 17220 128072 17276
rect 128120 17220 128176 17276
rect 128224 17220 128280 17276
rect 158736 17220 158792 17276
rect 158840 17220 158896 17276
rect 158944 17220 159000 17276
rect 189456 17220 189512 17276
rect 189560 17220 189616 17276
rect 189664 17220 189720 17276
rect 77308 17052 77364 17108
rect 78876 17052 78932 17108
rect 154812 16828 154868 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 127356 16436 127412 16492
rect 127460 16436 127516 16492
rect 127564 16436 127620 16492
rect 158076 16436 158132 16492
rect 158180 16436 158236 16492
rect 158284 16436 158340 16492
rect 188796 16436 188852 16492
rect 188900 16436 188956 16492
rect 189004 16436 189060 16492
rect 5136 15652 5192 15708
rect 5240 15652 5296 15708
rect 5344 15652 5400 15708
rect 35856 15652 35912 15708
rect 35960 15652 36016 15708
rect 36064 15652 36120 15708
rect 66576 15652 66632 15708
rect 66680 15652 66736 15708
rect 66784 15652 66840 15708
rect 97296 15652 97352 15708
rect 97400 15652 97456 15708
rect 97504 15652 97560 15708
rect 128016 15652 128072 15708
rect 128120 15652 128176 15708
rect 128224 15652 128280 15708
rect 158736 15652 158792 15708
rect 158840 15652 158896 15708
rect 158944 15652 159000 15708
rect 189456 15652 189512 15708
rect 189560 15652 189616 15708
rect 189664 15652 189720 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 127356 14868 127412 14924
rect 127460 14868 127516 14924
rect 127564 14868 127620 14924
rect 158076 14868 158132 14924
rect 158180 14868 158236 14924
rect 158284 14868 158340 14924
rect 188796 14868 188852 14924
rect 188900 14868 188956 14924
rect 189004 14868 189060 14924
rect 5136 14084 5192 14140
rect 5240 14084 5296 14140
rect 5344 14084 5400 14140
rect 35856 14084 35912 14140
rect 35960 14084 36016 14140
rect 36064 14084 36120 14140
rect 66576 14084 66632 14140
rect 66680 14084 66736 14140
rect 66784 14084 66840 14140
rect 97296 14084 97352 14140
rect 97400 14084 97456 14140
rect 97504 14084 97560 14140
rect 128016 14084 128072 14140
rect 128120 14084 128176 14140
rect 128224 14084 128280 14140
rect 158736 14084 158792 14140
rect 158840 14084 158896 14140
rect 158944 14084 159000 14140
rect 189456 14084 189512 14140
rect 189560 14084 189616 14140
rect 189664 14084 189720 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 127356 13300 127412 13356
rect 127460 13300 127516 13356
rect 127564 13300 127620 13356
rect 158076 13300 158132 13356
rect 158180 13300 158236 13356
rect 158284 13300 158340 13356
rect 188796 13300 188852 13356
rect 188900 13300 188956 13356
rect 189004 13300 189060 13356
rect 5136 12516 5192 12572
rect 5240 12516 5296 12572
rect 5344 12516 5400 12572
rect 35856 12516 35912 12572
rect 35960 12516 36016 12572
rect 36064 12516 36120 12572
rect 66576 12516 66632 12572
rect 66680 12516 66736 12572
rect 66784 12516 66840 12572
rect 97296 12516 97352 12572
rect 97400 12516 97456 12572
rect 97504 12516 97560 12572
rect 128016 12516 128072 12572
rect 128120 12516 128176 12572
rect 128224 12516 128280 12572
rect 158736 12516 158792 12572
rect 158840 12516 158896 12572
rect 158944 12516 159000 12572
rect 189456 12516 189512 12572
rect 189560 12516 189616 12572
rect 189664 12516 189720 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 127356 11732 127412 11788
rect 127460 11732 127516 11788
rect 127564 11732 127620 11788
rect 158076 11732 158132 11788
rect 158180 11732 158236 11788
rect 158284 11732 158340 11788
rect 188796 11732 188852 11788
rect 188900 11732 188956 11788
rect 189004 11732 189060 11788
rect 5136 10948 5192 11004
rect 5240 10948 5296 11004
rect 5344 10948 5400 11004
rect 35856 10948 35912 11004
rect 35960 10948 36016 11004
rect 36064 10948 36120 11004
rect 66576 10948 66632 11004
rect 66680 10948 66736 11004
rect 66784 10948 66840 11004
rect 97296 10948 97352 11004
rect 97400 10948 97456 11004
rect 97504 10948 97560 11004
rect 128016 10948 128072 11004
rect 128120 10948 128176 11004
rect 128224 10948 128280 11004
rect 158736 10948 158792 11004
rect 158840 10948 158896 11004
rect 158944 10948 159000 11004
rect 189456 10948 189512 11004
rect 189560 10948 189616 11004
rect 189664 10948 189720 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 127356 10164 127412 10220
rect 127460 10164 127516 10220
rect 127564 10164 127620 10220
rect 158076 10164 158132 10220
rect 158180 10164 158236 10220
rect 158284 10164 158340 10220
rect 188796 10164 188852 10220
rect 188900 10164 188956 10220
rect 189004 10164 189060 10220
rect 5136 9380 5192 9436
rect 5240 9380 5296 9436
rect 5344 9380 5400 9436
rect 35856 9380 35912 9436
rect 35960 9380 36016 9436
rect 36064 9380 36120 9436
rect 66576 9380 66632 9436
rect 66680 9380 66736 9436
rect 66784 9380 66840 9436
rect 97296 9380 97352 9436
rect 97400 9380 97456 9436
rect 97504 9380 97560 9436
rect 128016 9380 128072 9436
rect 128120 9380 128176 9436
rect 128224 9380 128280 9436
rect 158736 9380 158792 9436
rect 158840 9380 158896 9436
rect 158944 9380 159000 9436
rect 189456 9380 189512 9436
rect 189560 9380 189616 9436
rect 189664 9380 189720 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 127356 8596 127412 8652
rect 127460 8596 127516 8652
rect 127564 8596 127620 8652
rect 158076 8596 158132 8652
rect 158180 8596 158236 8652
rect 158284 8596 158340 8652
rect 188796 8596 188852 8652
rect 188900 8596 188956 8652
rect 189004 8596 189060 8652
rect 5136 7812 5192 7868
rect 5240 7812 5296 7868
rect 5344 7812 5400 7868
rect 35856 7812 35912 7868
rect 35960 7812 36016 7868
rect 36064 7812 36120 7868
rect 66576 7812 66632 7868
rect 66680 7812 66736 7868
rect 66784 7812 66840 7868
rect 97296 7812 97352 7868
rect 97400 7812 97456 7868
rect 97504 7812 97560 7868
rect 128016 7812 128072 7868
rect 128120 7812 128176 7868
rect 128224 7812 128280 7868
rect 158736 7812 158792 7868
rect 158840 7812 158896 7868
rect 158944 7812 159000 7868
rect 189456 7812 189512 7868
rect 189560 7812 189616 7868
rect 189664 7812 189720 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 127356 7028 127412 7084
rect 127460 7028 127516 7084
rect 127564 7028 127620 7084
rect 158076 7028 158132 7084
rect 158180 7028 158236 7084
rect 158284 7028 158340 7084
rect 188796 7028 188852 7084
rect 188900 7028 188956 7084
rect 189004 7028 189060 7084
rect 5136 6244 5192 6300
rect 5240 6244 5296 6300
rect 5344 6244 5400 6300
rect 35856 6244 35912 6300
rect 35960 6244 36016 6300
rect 36064 6244 36120 6300
rect 66576 6244 66632 6300
rect 66680 6244 66736 6300
rect 66784 6244 66840 6300
rect 97296 6244 97352 6300
rect 97400 6244 97456 6300
rect 97504 6244 97560 6300
rect 128016 6244 128072 6300
rect 128120 6244 128176 6300
rect 128224 6244 128280 6300
rect 158736 6244 158792 6300
rect 158840 6244 158896 6300
rect 158944 6244 159000 6300
rect 189456 6244 189512 6300
rect 189560 6244 189616 6300
rect 189664 6244 189720 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 127356 5460 127412 5516
rect 127460 5460 127516 5516
rect 127564 5460 127620 5516
rect 158076 5460 158132 5516
rect 158180 5460 158236 5516
rect 158284 5460 158340 5516
rect 188796 5460 188852 5516
rect 188900 5460 188956 5516
rect 189004 5460 189060 5516
rect 5136 4676 5192 4732
rect 5240 4676 5296 4732
rect 5344 4676 5400 4732
rect 35856 4676 35912 4732
rect 35960 4676 36016 4732
rect 36064 4676 36120 4732
rect 66576 4676 66632 4732
rect 66680 4676 66736 4732
rect 66784 4676 66840 4732
rect 97296 4676 97352 4732
rect 97400 4676 97456 4732
rect 97504 4676 97560 4732
rect 128016 4676 128072 4732
rect 128120 4676 128176 4732
rect 128224 4676 128280 4732
rect 158736 4676 158792 4732
rect 158840 4676 158896 4732
rect 158944 4676 159000 4732
rect 189456 4676 189512 4732
rect 189560 4676 189616 4732
rect 189664 4676 189720 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 127356 3892 127412 3948
rect 127460 3892 127516 3948
rect 127564 3892 127620 3948
rect 158076 3892 158132 3948
rect 158180 3892 158236 3948
rect 158284 3892 158340 3948
rect 188796 3892 188852 3948
rect 188900 3892 188956 3948
rect 189004 3892 189060 3948
rect 5136 3108 5192 3164
rect 5240 3108 5296 3164
rect 5344 3108 5400 3164
rect 35856 3108 35912 3164
rect 35960 3108 36016 3164
rect 36064 3108 36120 3164
rect 66576 3108 66632 3164
rect 66680 3108 66736 3164
rect 66784 3108 66840 3164
rect 97296 3108 97352 3164
rect 97400 3108 97456 3164
rect 97504 3108 97560 3164
rect 128016 3108 128072 3164
rect 128120 3108 128176 3164
rect 128224 3108 128280 3164
rect 158736 3108 158792 3164
rect 158840 3108 158896 3164
rect 158944 3108 159000 3164
rect 189456 3108 189512 3164
rect 189560 3108 189616 3164
rect 189664 3108 189720 3164
<< metal4 >>
rect 4448 156044 4768 156860
rect 4448 155988 4476 156044
rect 4532 155988 4580 156044
rect 4636 155988 4684 156044
rect 4740 155988 4768 156044
rect 4448 154476 4768 155988
rect 4448 154420 4476 154476
rect 4532 154420 4580 154476
rect 4636 154420 4684 154476
rect 4740 154420 4768 154476
rect 4448 152908 4768 154420
rect 4448 152852 4476 152908
rect 4532 152852 4580 152908
rect 4636 152852 4684 152908
rect 4740 152852 4768 152908
rect 4448 151340 4768 152852
rect 4448 151284 4476 151340
rect 4532 151284 4580 151340
rect 4636 151284 4684 151340
rect 4740 151284 4768 151340
rect 4448 149772 4768 151284
rect 4448 149716 4476 149772
rect 4532 149716 4580 149772
rect 4636 149716 4684 149772
rect 4740 149716 4768 149772
rect 4448 148204 4768 149716
rect 4448 148148 4476 148204
rect 4532 148148 4580 148204
rect 4636 148148 4684 148204
rect 4740 148148 4768 148204
rect 4448 146636 4768 148148
rect 4448 146580 4476 146636
rect 4532 146580 4580 146636
rect 4636 146580 4684 146636
rect 4740 146580 4768 146636
rect 4448 145068 4768 146580
rect 4448 145012 4476 145068
rect 4532 145012 4580 145068
rect 4636 145012 4684 145068
rect 4740 145012 4768 145068
rect 4448 143500 4768 145012
rect 4448 143444 4476 143500
rect 4532 143444 4580 143500
rect 4636 143444 4684 143500
rect 4740 143444 4768 143500
rect 4448 141932 4768 143444
rect 4448 141876 4476 141932
rect 4532 141876 4580 141932
rect 4636 141876 4684 141932
rect 4740 141876 4768 141932
rect 4448 140364 4768 141876
rect 4448 140308 4476 140364
rect 4532 140308 4580 140364
rect 4636 140308 4684 140364
rect 4740 140308 4768 140364
rect 4448 138796 4768 140308
rect 4448 138740 4476 138796
rect 4532 138740 4580 138796
rect 4636 138740 4684 138796
rect 4740 138740 4768 138796
rect 4448 137228 4768 138740
rect 4448 137172 4476 137228
rect 4532 137172 4580 137228
rect 4636 137172 4684 137228
rect 4740 137172 4768 137228
rect 4448 135660 4768 137172
rect 4448 135604 4476 135660
rect 4532 135604 4580 135660
rect 4636 135604 4684 135660
rect 4740 135604 4768 135660
rect 4448 134092 4768 135604
rect 4448 134036 4476 134092
rect 4532 134036 4580 134092
rect 4636 134036 4684 134092
rect 4740 134036 4768 134092
rect 4448 132524 4768 134036
rect 4448 132468 4476 132524
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4740 132468 4768 132524
rect 4448 130956 4768 132468
rect 4448 130900 4476 130956
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4740 130900 4768 130956
rect 4448 129388 4768 130900
rect 4448 129332 4476 129388
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4740 129332 4768 129388
rect 4448 129142 4768 129332
rect 4448 129086 4476 129142
rect 4532 129086 4580 129142
rect 4636 129086 4684 129142
rect 4740 129086 4768 129142
rect 4448 129038 4768 129086
rect 4448 128982 4476 129038
rect 4532 128982 4580 129038
rect 4636 128982 4684 129038
rect 4740 128982 4768 129038
rect 4448 128934 4768 128982
rect 4448 128878 4476 128934
rect 4532 128878 4580 128934
rect 4636 128878 4684 128934
rect 4740 128878 4768 128934
rect 4448 127820 4768 128878
rect 4448 127764 4476 127820
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4740 127764 4768 127820
rect 4448 126252 4768 127764
rect 4448 126196 4476 126252
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4740 126196 4768 126252
rect 4448 124684 4768 126196
rect 4448 124628 4476 124684
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4740 124628 4768 124684
rect 4448 123116 4768 124628
rect 4448 123060 4476 123116
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4740 123060 4768 123116
rect 4448 121548 4768 123060
rect 4448 121492 4476 121548
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4740 121492 4768 121548
rect 4448 119980 4768 121492
rect 4448 119924 4476 119980
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4740 119924 4768 119980
rect 4448 118412 4768 119924
rect 4448 118356 4476 118412
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4740 118356 4768 118412
rect 4448 116844 4768 118356
rect 4448 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4768 116844
rect 4448 115276 4768 116788
rect 4448 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4768 115276
rect 4448 113708 4768 115220
rect 4448 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4768 113708
rect 4448 112140 4768 113652
rect 4448 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4768 112140
rect 4448 110572 4768 112084
rect 4448 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4768 110572
rect 4448 109004 4768 110516
rect 4448 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4768 109004
rect 4448 107436 4768 108948
rect 4448 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4768 107436
rect 4448 105868 4768 107380
rect 4448 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4768 105868
rect 4448 104300 4768 105812
rect 4448 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4768 104300
rect 4448 102732 4768 104244
rect 4448 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4768 102732
rect 4448 101164 4768 102676
rect 4448 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4768 101164
rect 4448 99596 4768 101108
rect 4448 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4768 99596
rect 4448 98506 4768 99540
rect 4448 98450 4476 98506
rect 4532 98450 4580 98506
rect 4636 98450 4684 98506
rect 4740 98450 4768 98506
rect 4448 98402 4768 98450
rect 4448 98346 4476 98402
rect 4532 98346 4580 98402
rect 4636 98346 4684 98402
rect 4740 98346 4768 98402
rect 4448 98298 4768 98346
rect 4448 98242 4476 98298
rect 4532 98242 4580 98298
rect 4636 98242 4684 98298
rect 4740 98242 4768 98298
rect 4448 98028 4768 98242
rect 4448 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4768 98028
rect 4448 96460 4768 97972
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 67870 4768 68180
rect 4448 67814 4476 67870
rect 4532 67814 4580 67870
rect 4636 67814 4684 67870
rect 4740 67814 4768 67870
rect 4448 67766 4768 67814
rect 4448 67710 4476 67766
rect 4532 67710 4580 67766
rect 4636 67710 4684 67766
rect 4740 67710 4768 67766
rect 4448 67662 4768 67710
rect 4448 67606 4476 67662
rect 4532 67606 4580 67662
rect 4636 67606 4684 67662
rect 4740 67606 4768 67662
rect 4448 66668 4768 67606
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 37234 4768 38388
rect 4448 37178 4476 37234
rect 4532 37178 4580 37234
rect 4636 37178 4684 37234
rect 4740 37178 4768 37234
rect 4448 37130 4768 37178
rect 4448 37074 4476 37130
rect 4532 37074 4580 37130
rect 4636 37074 4684 37130
rect 4740 37074 4768 37130
rect 4448 37026 4768 37074
rect 4448 36970 4476 37026
rect 4532 36970 4580 37026
rect 4636 36970 4684 37026
rect 4740 36970 4768 37026
rect 4448 36876 4768 36970
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 6598 4768 7028
rect 4448 6542 4476 6598
rect 4532 6542 4580 6598
rect 4636 6542 4684 6598
rect 4740 6542 4768 6598
rect 4448 6494 4768 6542
rect 4448 6438 4476 6494
rect 4532 6438 4580 6494
rect 4636 6438 4684 6494
rect 4740 6438 4768 6494
rect 4448 6390 4768 6438
rect 4448 6334 4476 6390
rect 4532 6334 4580 6390
rect 4636 6334 4684 6390
rect 4740 6334 4768 6390
rect 4448 5516 4768 6334
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 5108 156828 5428 156860
rect 5108 156772 5136 156828
rect 5192 156772 5240 156828
rect 5296 156772 5344 156828
rect 5400 156772 5428 156828
rect 5108 155260 5428 156772
rect 5108 155204 5136 155260
rect 5192 155204 5240 155260
rect 5296 155204 5344 155260
rect 5400 155204 5428 155260
rect 5108 153692 5428 155204
rect 5108 153636 5136 153692
rect 5192 153636 5240 153692
rect 5296 153636 5344 153692
rect 5400 153636 5428 153692
rect 5108 152124 5428 153636
rect 5108 152068 5136 152124
rect 5192 152068 5240 152124
rect 5296 152068 5344 152124
rect 5400 152068 5428 152124
rect 5108 150556 5428 152068
rect 5108 150500 5136 150556
rect 5192 150500 5240 150556
rect 5296 150500 5344 150556
rect 5400 150500 5428 150556
rect 5108 148988 5428 150500
rect 5108 148932 5136 148988
rect 5192 148932 5240 148988
rect 5296 148932 5344 148988
rect 5400 148932 5428 148988
rect 5108 147420 5428 148932
rect 5108 147364 5136 147420
rect 5192 147364 5240 147420
rect 5296 147364 5344 147420
rect 5400 147364 5428 147420
rect 5108 145852 5428 147364
rect 5108 145796 5136 145852
rect 5192 145796 5240 145852
rect 5296 145796 5344 145852
rect 5400 145796 5428 145852
rect 5108 144284 5428 145796
rect 5108 144228 5136 144284
rect 5192 144228 5240 144284
rect 5296 144228 5344 144284
rect 5400 144228 5428 144284
rect 5108 142716 5428 144228
rect 5108 142660 5136 142716
rect 5192 142660 5240 142716
rect 5296 142660 5344 142716
rect 5400 142660 5428 142716
rect 5108 141148 5428 142660
rect 5108 141092 5136 141148
rect 5192 141092 5240 141148
rect 5296 141092 5344 141148
rect 5400 141092 5428 141148
rect 5108 139580 5428 141092
rect 5108 139524 5136 139580
rect 5192 139524 5240 139580
rect 5296 139524 5344 139580
rect 5400 139524 5428 139580
rect 5108 138012 5428 139524
rect 5108 137956 5136 138012
rect 5192 137956 5240 138012
rect 5296 137956 5344 138012
rect 5400 137956 5428 138012
rect 5108 136444 5428 137956
rect 5108 136388 5136 136444
rect 5192 136388 5240 136444
rect 5296 136388 5344 136444
rect 5400 136388 5428 136444
rect 5108 134876 5428 136388
rect 5108 134820 5136 134876
rect 5192 134820 5240 134876
rect 5296 134820 5344 134876
rect 5400 134820 5428 134876
rect 5108 133308 5428 134820
rect 5108 133252 5136 133308
rect 5192 133252 5240 133308
rect 5296 133252 5344 133308
rect 5400 133252 5428 133308
rect 5108 131740 5428 133252
rect 5108 131684 5136 131740
rect 5192 131684 5240 131740
rect 5296 131684 5344 131740
rect 5400 131684 5428 131740
rect 5108 130172 5428 131684
rect 5108 130116 5136 130172
rect 5192 130116 5240 130172
rect 5296 130116 5344 130172
rect 5400 130116 5428 130172
rect 5108 129802 5428 130116
rect 35168 156044 35488 156860
rect 35168 155988 35196 156044
rect 35252 155988 35300 156044
rect 35356 155988 35404 156044
rect 35460 155988 35488 156044
rect 35168 154476 35488 155988
rect 35168 154420 35196 154476
rect 35252 154420 35300 154476
rect 35356 154420 35404 154476
rect 35460 154420 35488 154476
rect 35168 152908 35488 154420
rect 35168 152852 35196 152908
rect 35252 152852 35300 152908
rect 35356 152852 35404 152908
rect 35460 152852 35488 152908
rect 35168 151340 35488 152852
rect 35168 151284 35196 151340
rect 35252 151284 35300 151340
rect 35356 151284 35404 151340
rect 35460 151284 35488 151340
rect 35168 149772 35488 151284
rect 35168 149716 35196 149772
rect 35252 149716 35300 149772
rect 35356 149716 35404 149772
rect 35460 149716 35488 149772
rect 35168 148204 35488 149716
rect 35168 148148 35196 148204
rect 35252 148148 35300 148204
rect 35356 148148 35404 148204
rect 35460 148148 35488 148204
rect 35168 146636 35488 148148
rect 35168 146580 35196 146636
rect 35252 146580 35300 146636
rect 35356 146580 35404 146636
rect 35460 146580 35488 146636
rect 35168 145068 35488 146580
rect 35168 145012 35196 145068
rect 35252 145012 35300 145068
rect 35356 145012 35404 145068
rect 35460 145012 35488 145068
rect 5108 129746 5136 129802
rect 5192 129746 5240 129802
rect 5296 129746 5344 129802
rect 5400 129746 5428 129802
rect 5108 129698 5428 129746
rect 5108 129642 5136 129698
rect 5192 129642 5240 129698
rect 5296 129642 5344 129698
rect 5400 129642 5428 129698
rect 5108 129594 5428 129642
rect 5108 129538 5136 129594
rect 5192 129538 5240 129594
rect 5296 129538 5344 129594
rect 5400 129538 5428 129594
rect 5108 128604 5428 129538
rect 20000 129802 20340 129830
rect 20000 129746 20038 129802
rect 20094 129746 20142 129802
rect 20198 129746 20246 129802
rect 20302 129746 20340 129802
rect 20000 129698 20340 129746
rect 20000 129642 20038 129698
rect 20094 129642 20142 129698
rect 20198 129642 20246 129698
rect 20302 129642 20340 129698
rect 20000 129594 20340 129642
rect 20000 129538 20038 129594
rect 20094 129538 20142 129594
rect 20198 129538 20246 129594
rect 20302 129538 20340 129594
rect 20000 129510 20340 129538
rect 20660 129142 21000 129170
rect 20660 129086 20698 129142
rect 20754 129086 20802 129142
rect 20858 129086 20906 129142
rect 20962 129086 21000 129142
rect 20660 129038 21000 129086
rect 20660 128982 20698 129038
rect 20754 128982 20802 129038
rect 20858 128982 20906 129038
rect 20962 128982 21000 129038
rect 20660 128934 21000 128982
rect 20660 128878 20698 128934
rect 20754 128878 20802 128934
rect 20858 128878 20906 128934
rect 20962 128878 21000 128934
rect 20660 128850 21000 128878
rect 35168 129142 35488 145012
rect 35168 129086 35196 129142
rect 35252 129086 35300 129142
rect 35356 129086 35404 129142
rect 35460 129086 35488 129142
rect 35168 129038 35488 129086
rect 35168 128982 35196 129038
rect 35252 128982 35300 129038
rect 35356 128982 35404 129038
rect 35460 128982 35488 129038
rect 35168 128934 35488 128982
rect 35168 128878 35196 128934
rect 35252 128878 35300 128934
rect 35356 128878 35404 128934
rect 35460 128878 35488 128934
rect 5108 128548 5136 128604
rect 5192 128548 5240 128604
rect 5296 128548 5344 128604
rect 5400 128548 5428 128604
rect 5108 127036 5428 128548
rect 5108 126980 5136 127036
rect 5192 126980 5240 127036
rect 5296 126980 5344 127036
rect 5400 126980 5428 127036
rect 5108 125468 5428 126980
rect 5108 125412 5136 125468
rect 5192 125412 5240 125468
rect 5296 125412 5344 125468
rect 5400 125412 5428 125468
rect 5108 123900 5428 125412
rect 5108 123844 5136 123900
rect 5192 123844 5240 123900
rect 5296 123844 5344 123900
rect 5400 123844 5428 123900
rect 5108 122332 5428 123844
rect 5108 122276 5136 122332
rect 5192 122276 5240 122332
rect 5296 122276 5344 122332
rect 5400 122276 5428 122332
rect 5108 120764 5428 122276
rect 5108 120708 5136 120764
rect 5192 120708 5240 120764
rect 5296 120708 5344 120764
rect 5400 120708 5428 120764
rect 5108 119196 5428 120708
rect 5108 119140 5136 119196
rect 5192 119140 5240 119196
rect 5296 119140 5344 119196
rect 5400 119140 5428 119196
rect 5108 117628 5428 119140
rect 5108 117572 5136 117628
rect 5192 117572 5240 117628
rect 5296 117572 5344 117628
rect 5400 117572 5428 117628
rect 5108 116060 5428 117572
rect 5108 116004 5136 116060
rect 5192 116004 5240 116060
rect 5296 116004 5344 116060
rect 5400 116004 5428 116060
rect 5108 114492 5428 116004
rect 5108 114436 5136 114492
rect 5192 114436 5240 114492
rect 5296 114436 5344 114492
rect 5400 114436 5428 114492
rect 5108 112924 5428 114436
rect 5108 112868 5136 112924
rect 5192 112868 5240 112924
rect 5296 112868 5344 112924
rect 5400 112868 5428 112924
rect 5108 111356 5428 112868
rect 5108 111300 5136 111356
rect 5192 111300 5240 111356
rect 5296 111300 5344 111356
rect 5400 111300 5428 111356
rect 5108 109788 5428 111300
rect 5108 109732 5136 109788
rect 5192 109732 5240 109788
rect 5296 109732 5344 109788
rect 5400 109732 5428 109788
rect 5108 108220 5428 109732
rect 5108 108164 5136 108220
rect 5192 108164 5240 108220
rect 5296 108164 5344 108220
rect 5400 108164 5428 108220
rect 5108 106652 5428 108164
rect 5108 106596 5136 106652
rect 5192 106596 5240 106652
rect 5296 106596 5344 106652
rect 5400 106596 5428 106652
rect 5108 105084 5428 106596
rect 5108 105028 5136 105084
rect 5192 105028 5240 105084
rect 5296 105028 5344 105084
rect 5400 105028 5428 105084
rect 5108 103516 5428 105028
rect 5108 103460 5136 103516
rect 5192 103460 5240 103516
rect 5296 103460 5344 103516
rect 5400 103460 5428 103516
rect 5108 101948 5428 103460
rect 5108 101892 5136 101948
rect 5192 101892 5240 101948
rect 5296 101892 5344 101948
rect 5400 101892 5428 101948
rect 5108 100380 5428 101892
rect 5108 100324 5136 100380
rect 5192 100324 5240 100380
rect 5296 100324 5344 100380
rect 5400 100324 5428 100380
rect 5108 99166 5428 100324
rect 5108 99110 5136 99166
rect 5192 99110 5240 99166
rect 5296 99110 5344 99166
rect 5400 99110 5428 99166
rect 5108 99062 5428 99110
rect 5108 99006 5136 99062
rect 5192 99006 5240 99062
rect 5296 99006 5344 99062
rect 5400 99006 5428 99062
rect 5108 98958 5428 99006
rect 5108 98902 5136 98958
rect 5192 98902 5240 98958
rect 5296 98902 5344 98958
rect 5400 98902 5428 98958
rect 5108 98812 5428 98902
rect 20000 99166 20340 99194
rect 20000 99110 20038 99166
rect 20094 99110 20142 99166
rect 20198 99110 20246 99166
rect 20302 99110 20340 99166
rect 20000 99062 20340 99110
rect 20000 99006 20038 99062
rect 20094 99006 20142 99062
rect 20198 99006 20246 99062
rect 20302 99006 20340 99062
rect 20000 98958 20340 99006
rect 20000 98902 20038 98958
rect 20094 98902 20142 98958
rect 20198 98902 20246 98958
rect 20302 98902 20340 98958
rect 20000 98874 20340 98902
rect 5108 98756 5136 98812
rect 5192 98756 5240 98812
rect 5296 98756 5344 98812
rect 5400 98756 5428 98812
rect 5108 97244 5428 98756
rect 20660 98506 21000 98534
rect 20660 98450 20698 98506
rect 20754 98450 20802 98506
rect 20858 98450 20906 98506
rect 20962 98450 21000 98506
rect 20660 98402 21000 98450
rect 20660 98346 20698 98402
rect 20754 98346 20802 98402
rect 20858 98346 20906 98402
rect 20962 98346 21000 98402
rect 20660 98298 21000 98346
rect 20660 98242 20698 98298
rect 20754 98242 20802 98298
rect 20858 98242 20906 98298
rect 20962 98242 21000 98298
rect 20660 98214 21000 98242
rect 35168 98506 35488 128878
rect 35168 98450 35196 98506
rect 35252 98450 35300 98506
rect 35356 98450 35404 98506
rect 35460 98450 35488 98506
rect 35168 98402 35488 98450
rect 35168 98346 35196 98402
rect 35252 98346 35300 98402
rect 35356 98346 35404 98402
rect 35460 98346 35488 98402
rect 35168 98298 35488 98346
rect 35168 98242 35196 98298
rect 35252 98242 35300 98298
rect 35356 98242 35404 98298
rect 35460 98242 35488 98298
rect 5108 97188 5136 97244
rect 5192 97188 5240 97244
rect 5296 97188 5344 97244
rect 5400 97188 5428 97244
rect 5108 95676 5428 97188
rect 5108 95620 5136 95676
rect 5192 95620 5240 95676
rect 5296 95620 5344 95676
rect 5400 95620 5428 95676
rect 5108 94108 5428 95620
rect 5108 94052 5136 94108
rect 5192 94052 5240 94108
rect 5296 94052 5344 94108
rect 5400 94052 5428 94108
rect 5108 92540 5428 94052
rect 5108 92484 5136 92540
rect 5192 92484 5240 92540
rect 5296 92484 5344 92540
rect 5400 92484 5428 92540
rect 5108 90972 5428 92484
rect 5108 90916 5136 90972
rect 5192 90916 5240 90972
rect 5296 90916 5344 90972
rect 5400 90916 5428 90972
rect 5108 89404 5428 90916
rect 5108 89348 5136 89404
rect 5192 89348 5240 89404
rect 5296 89348 5344 89404
rect 5400 89348 5428 89404
rect 5108 87836 5428 89348
rect 5108 87780 5136 87836
rect 5192 87780 5240 87836
rect 5296 87780 5344 87836
rect 5400 87780 5428 87836
rect 5108 86268 5428 87780
rect 5108 86212 5136 86268
rect 5192 86212 5240 86268
rect 5296 86212 5344 86268
rect 5400 86212 5428 86268
rect 5108 84700 5428 86212
rect 5108 84644 5136 84700
rect 5192 84644 5240 84700
rect 5296 84644 5344 84700
rect 5400 84644 5428 84700
rect 5108 83132 5428 84644
rect 5108 83076 5136 83132
rect 5192 83076 5240 83132
rect 5296 83076 5344 83132
rect 5400 83076 5428 83132
rect 5108 81564 5428 83076
rect 5108 81508 5136 81564
rect 5192 81508 5240 81564
rect 5296 81508 5344 81564
rect 5400 81508 5428 81564
rect 5108 79996 5428 81508
rect 5108 79940 5136 79996
rect 5192 79940 5240 79996
rect 5296 79940 5344 79996
rect 5400 79940 5428 79996
rect 5108 78428 5428 79940
rect 5108 78372 5136 78428
rect 5192 78372 5240 78428
rect 5296 78372 5344 78428
rect 5400 78372 5428 78428
rect 5108 76860 5428 78372
rect 5108 76804 5136 76860
rect 5192 76804 5240 76860
rect 5296 76804 5344 76860
rect 5400 76804 5428 76860
rect 5108 75292 5428 76804
rect 5108 75236 5136 75292
rect 5192 75236 5240 75292
rect 5296 75236 5344 75292
rect 5400 75236 5428 75292
rect 5108 73724 5428 75236
rect 5108 73668 5136 73724
rect 5192 73668 5240 73724
rect 5296 73668 5344 73724
rect 5400 73668 5428 73724
rect 5108 72156 5428 73668
rect 5108 72100 5136 72156
rect 5192 72100 5240 72156
rect 5296 72100 5344 72156
rect 5400 72100 5428 72156
rect 5108 70588 5428 72100
rect 5108 70532 5136 70588
rect 5192 70532 5240 70588
rect 5296 70532 5344 70588
rect 5400 70532 5428 70588
rect 5108 69020 5428 70532
rect 5108 68964 5136 69020
rect 5192 68964 5240 69020
rect 5296 68964 5344 69020
rect 5400 68964 5428 69020
rect 5108 68530 5428 68964
rect 5108 68474 5136 68530
rect 5192 68474 5240 68530
rect 5296 68474 5344 68530
rect 5400 68474 5428 68530
rect 5108 68426 5428 68474
rect 5108 68370 5136 68426
rect 5192 68370 5240 68426
rect 5296 68370 5344 68426
rect 5400 68370 5428 68426
rect 5108 68322 5428 68370
rect 5108 68266 5136 68322
rect 5192 68266 5240 68322
rect 5296 68266 5344 68322
rect 5400 68266 5428 68322
rect 5108 67452 5428 68266
rect 20000 68530 20340 68558
rect 20000 68474 20038 68530
rect 20094 68474 20142 68530
rect 20198 68474 20246 68530
rect 20302 68474 20340 68530
rect 20000 68426 20340 68474
rect 20000 68370 20038 68426
rect 20094 68370 20142 68426
rect 20198 68370 20246 68426
rect 20302 68370 20340 68426
rect 20000 68322 20340 68370
rect 20000 68266 20038 68322
rect 20094 68266 20142 68322
rect 20198 68266 20246 68322
rect 20302 68266 20340 68322
rect 20000 68238 20340 68266
rect 20660 67870 21000 67898
rect 20660 67814 20698 67870
rect 20754 67814 20802 67870
rect 20858 67814 20906 67870
rect 20962 67814 21000 67870
rect 20660 67766 21000 67814
rect 20660 67710 20698 67766
rect 20754 67710 20802 67766
rect 20858 67710 20906 67766
rect 20962 67710 21000 67766
rect 20660 67662 21000 67710
rect 20660 67606 20698 67662
rect 20754 67606 20802 67662
rect 20858 67606 20906 67662
rect 20962 67606 21000 67662
rect 20660 67578 21000 67606
rect 35168 67870 35488 98242
rect 35168 67814 35196 67870
rect 35252 67814 35300 67870
rect 35356 67814 35404 67870
rect 35460 67814 35488 67870
rect 35168 67766 35488 67814
rect 35168 67710 35196 67766
rect 35252 67710 35300 67766
rect 35356 67710 35404 67766
rect 35460 67710 35488 67766
rect 35168 67662 35488 67710
rect 35168 67606 35196 67662
rect 35252 67606 35300 67662
rect 35356 67606 35404 67662
rect 35460 67606 35488 67662
rect 5108 67396 5136 67452
rect 5192 67396 5240 67452
rect 5296 67396 5344 67452
rect 5400 67396 5428 67452
rect 5108 65884 5428 67396
rect 5108 65828 5136 65884
rect 5192 65828 5240 65884
rect 5296 65828 5344 65884
rect 5400 65828 5428 65884
rect 5108 64316 5428 65828
rect 5108 64260 5136 64316
rect 5192 64260 5240 64316
rect 5296 64260 5344 64316
rect 5400 64260 5428 64316
rect 5108 62748 5428 64260
rect 5108 62692 5136 62748
rect 5192 62692 5240 62748
rect 5296 62692 5344 62748
rect 5400 62692 5428 62748
rect 5108 61180 5428 62692
rect 5108 61124 5136 61180
rect 5192 61124 5240 61180
rect 5296 61124 5344 61180
rect 5400 61124 5428 61180
rect 5108 59612 5428 61124
rect 5108 59556 5136 59612
rect 5192 59556 5240 59612
rect 5296 59556 5344 59612
rect 5400 59556 5428 59612
rect 5108 58044 5428 59556
rect 5108 57988 5136 58044
rect 5192 57988 5240 58044
rect 5296 57988 5344 58044
rect 5400 57988 5428 58044
rect 5108 56476 5428 57988
rect 5108 56420 5136 56476
rect 5192 56420 5240 56476
rect 5296 56420 5344 56476
rect 5400 56420 5428 56476
rect 5108 54908 5428 56420
rect 5108 54852 5136 54908
rect 5192 54852 5240 54908
rect 5296 54852 5344 54908
rect 5400 54852 5428 54908
rect 5108 53340 5428 54852
rect 5108 53284 5136 53340
rect 5192 53284 5240 53340
rect 5296 53284 5344 53340
rect 5400 53284 5428 53340
rect 5108 51772 5428 53284
rect 5108 51716 5136 51772
rect 5192 51716 5240 51772
rect 5296 51716 5344 51772
rect 5400 51716 5428 51772
rect 5108 50204 5428 51716
rect 5108 50148 5136 50204
rect 5192 50148 5240 50204
rect 5296 50148 5344 50204
rect 5400 50148 5428 50204
rect 5108 48636 5428 50148
rect 5108 48580 5136 48636
rect 5192 48580 5240 48636
rect 5296 48580 5344 48636
rect 5400 48580 5428 48636
rect 5108 47068 5428 48580
rect 5108 47012 5136 47068
rect 5192 47012 5240 47068
rect 5296 47012 5344 47068
rect 5400 47012 5428 47068
rect 5108 45500 5428 47012
rect 5108 45444 5136 45500
rect 5192 45444 5240 45500
rect 5296 45444 5344 45500
rect 5400 45444 5428 45500
rect 5108 43932 5428 45444
rect 5108 43876 5136 43932
rect 5192 43876 5240 43932
rect 5296 43876 5344 43932
rect 5400 43876 5428 43932
rect 5108 42364 5428 43876
rect 5108 42308 5136 42364
rect 5192 42308 5240 42364
rect 5296 42308 5344 42364
rect 5400 42308 5428 42364
rect 5108 40796 5428 42308
rect 5108 40740 5136 40796
rect 5192 40740 5240 40796
rect 5296 40740 5344 40796
rect 5400 40740 5428 40796
rect 5108 39228 5428 40740
rect 5108 39172 5136 39228
rect 5192 39172 5240 39228
rect 5296 39172 5344 39228
rect 5400 39172 5428 39228
rect 5108 37894 5428 39172
rect 5108 37838 5136 37894
rect 5192 37838 5240 37894
rect 5296 37838 5344 37894
rect 5400 37838 5428 37894
rect 5108 37790 5428 37838
rect 5108 37734 5136 37790
rect 5192 37734 5240 37790
rect 5296 37734 5344 37790
rect 5400 37734 5428 37790
rect 5108 37686 5428 37734
rect 5108 37604 5136 37686
rect 5192 37604 5240 37686
rect 5296 37604 5344 37686
rect 5400 37604 5428 37686
rect 5108 36092 5428 37604
rect 20000 37894 20340 37922
rect 20000 37838 20038 37894
rect 20094 37838 20142 37894
rect 20198 37838 20246 37894
rect 20302 37838 20340 37894
rect 20000 37790 20340 37838
rect 20000 37734 20038 37790
rect 20094 37734 20142 37790
rect 20198 37734 20246 37790
rect 20302 37734 20340 37790
rect 20000 37686 20340 37734
rect 20000 37630 20038 37686
rect 20094 37630 20142 37686
rect 20198 37630 20246 37686
rect 20302 37630 20340 37686
rect 20000 37602 20340 37630
rect 29052 37894 29128 37922
rect 29052 37838 29062 37894
rect 29118 37838 29128 37894
rect 29052 37790 29128 37838
rect 29052 37734 29062 37790
rect 29118 37734 29128 37790
rect 29052 37686 29128 37734
rect 29052 37630 29062 37686
rect 29118 37630 29128 37686
rect 29052 37602 29128 37630
rect 20660 37234 21000 37262
rect 20660 37178 20698 37234
rect 20754 37178 20802 37234
rect 20858 37178 20906 37234
rect 20962 37178 21000 37234
rect 20660 37130 21000 37178
rect 20660 37074 20698 37130
rect 20754 37074 20802 37130
rect 20858 37074 20906 37130
rect 20962 37074 21000 37130
rect 20660 37026 21000 37074
rect 20660 36970 20698 37026
rect 20754 36970 20802 37026
rect 20858 36970 20906 37026
rect 20962 36970 21000 37026
rect 20660 36942 21000 36970
rect 35168 37234 35488 67606
rect 35168 37178 35196 37234
rect 35252 37178 35300 37234
rect 35356 37178 35404 37234
rect 35460 37178 35488 37234
rect 35168 37130 35488 37178
rect 35168 37074 35196 37130
rect 35252 37074 35300 37130
rect 35356 37074 35404 37130
rect 35460 37074 35488 37130
rect 35168 37026 35488 37074
rect 35168 36970 35196 37026
rect 35252 36970 35300 37026
rect 35356 36970 35404 37026
rect 35460 36970 35488 37026
rect 5108 36036 5136 36092
rect 5192 36036 5240 36092
rect 5296 36036 5344 36092
rect 5400 36036 5428 36092
rect 5108 34524 5428 36036
rect 5108 34468 5136 34524
rect 5192 34468 5240 34524
rect 5296 34468 5344 34524
rect 5400 34468 5428 34524
rect 5108 32956 5428 34468
rect 5108 32900 5136 32956
rect 5192 32900 5240 32956
rect 5296 32900 5344 32956
rect 5400 32900 5428 32956
rect 5108 31388 5428 32900
rect 5108 31332 5136 31388
rect 5192 31332 5240 31388
rect 5296 31332 5344 31388
rect 5400 31332 5428 31388
rect 5108 29820 5428 31332
rect 5108 29764 5136 29820
rect 5192 29764 5240 29820
rect 5296 29764 5344 29820
rect 5400 29764 5428 29820
rect 5108 28252 5428 29764
rect 5108 28196 5136 28252
rect 5192 28196 5240 28252
rect 5296 28196 5344 28252
rect 5400 28196 5428 28252
rect 5108 26684 5428 28196
rect 5108 26628 5136 26684
rect 5192 26628 5240 26684
rect 5296 26628 5344 26684
rect 5400 26628 5428 26684
rect 5108 25116 5428 26628
rect 5108 25060 5136 25116
rect 5192 25060 5240 25116
rect 5296 25060 5344 25116
rect 5400 25060 5428 25116
rect 5108 23548 5428 25060
rect 5108 23492 5136 23548
rect 5192 23492 5240 23548
rect 5296 23492 5344 23548
rect 5400 23492 5428 23548
rect 5108 21980 5428 23492
rect 5108 21924 5136 21980
rect 5192 21924 5240 21980
rect 5296 21924 5344 21980
rect 5400 21924 5428 21980
rect 5108 20412 5428 21924
rect 5108 20356 5136 20412
rect 5192 20356 5240 20412
rect 5296 20356 5344 20412
rect 5400 20356 5428 20412
rect 5108 18844 5428 20356
rect 5108 18788 5136 18844
rect 5192 18788 5240 18844
rect 5296 18788 5344 18844
rect 5400 18788 5428 18844
rect 5108 17276 5428 18788
rect 5108 17220 5136 17276
rect 5192 17220 5240 17276
rect 5296 17220 5344 17276
rect 5400 17220 5428 17276
rect 5108 15708 5428 17220
rect 5108 15652 5136 15708
rect 5192 15652 5240 15708
rect 5296 15652 5344 15708
rect 5400 15652 5428 15708
rect 5108 14140 5428 15652
rect 5108 14084 5136 14140
rect 5192 14084 5240 14140
rect 5296 14084 5344 14140
rect 5400 14084 5428 14140
rect 5108 12572 5428 14084
rect 5108 12516 5136 12572
rect 5192 12516 5240 12572
rect 5296 12516 5344 12572
rect 5400 12516 5428 12572
rect 5108 11004 5428 12516
rect 5108 10948 5136 11004
rect 5192 10948 5240 11004
rect 5296 10948 5344 11004
rect 5400 10948 5428 11004
rect 5108 9436 5428 10948
rect 5108 9380 5136 9436
rect 5192 9380 5240 9436
rect 5296 9380 5344 9436
rect 5400 9380 5428 9436
rect 5108 7868 5428 9380
rect 5108 7812 5136 7868
rect 5192 7812 5240 7868
rect 5296 7812 5344 7868
rect 5400 7812 5428 7868
rect 5108 7258 5428 7812
rect 5108 7202 5136 7258
rect 5192 7202 5240 7258
rect 5296 7202 5344 7258
rect 5400 7202 5428 7258
rect 5108 7154 5428 7202
rect 5108 7098 5136 7154
rect 5192 7098 5240 7154
rect 5296 7098 5344 7154
rect 5400 7098 5428 7154
rect 5108 7050 5428 7098
rect 5108 6994 5136 7050
rect 5192 6994 5240 7050
rect 5296 6994 5344 7050
rect 5400 6994 5428 7050
rect 5108 6300 5428 6994
rect 5108 6244 5136 6300
rect 5192 6244 5240 6300
rect 5296 6244 5344 6300
rect 5400 6244 5428 6300
rect 5108 4732 5428 6244
rect 5108 4676 5136 4732
rect 5192 4676 5240 4732
rect 5296 4676 5344 4732
rect 5400 4676 5428 4732
rect 5108 3164 5428 4676
rect 5108 3108 5136 3164
rect 5192 3108 5240 3164
rect 5296 3108 5344 3164
rect 5400 3108 5428 3164
rect 5108 3076 5428 3108
rect 35168 16492 35488 36970
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 6598 35488 7028
rect 35168 6542 35196 6598
rect 35252 6542 35300 6598
rect 35356 6542 35404 6598
rect 35460 6542 35488 6598
rect 35168 6494 35488 6542
rect 35168 6438 35196 6494
rect 35252 6438 35300 6494
rect 35356 6438 35404 6494
rect 35460 6438 35488 6494
rect 35168 6390 35488 6438
rect 35168 6334 35196 6390
rect 35252 6334 35300 6390
rect 35356 6334 35404 6390
rect 35460 6334 35488 6390
rect 35168 5516 35488 6334
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 35828 156828 36148 156860
rect 35828 156772 35856 156828
rect 35912 156772 35960 156828
rect 36016 156772 36064 156828
rect 36120 156772 36148 156828
rect 35828 155260 36148 156772
rect 35828 155204 35856 155260
rect 35912 155204 35960 155260
rect 36016 155204 36064 155260
rect 36120 155204 36148 155260
rect 35828 153692 36148 155204
rect 35828 153636 35856 153692
rect 35912 153636 35960 153692
rect 36016 153636 36064 153692
rect 36120 153636 36148 153692
rect 35828 152124 36148 153636
rect 35828 152068 35856 152124
rect 35912 152068 35960 152124
rect 36016 152068 36064 152124
rect 36120 152068 36148 152124
rect 35828 150556 36148 152068
rect 35828 150500 35856 150556
rect 35912 150500 35960 150556
rect 36016 150500 36064 150556
rect 36120 150500 36148 150556
rect 35828 148988 36148 150500
rect 35828 148932 35856 148988
rect 35912 148932 35960 148988
rect 36016 148932 36064 148988
rect 36120 148932 36148 148988
rect 35828 147420 36148 148932
rect 35828 147364 35856 147420
rect 35912 147364 35960 147420
rect 36016 147364 36064 147420
rect 36120 147364 36148 147420
rect 35828 145852 36148 147364
rect 35828 145796 35856 145852
rect 35912 145796 35960 145852
rect 36016 145796 36064 145852
rect 36120 145796 36148 145852
rect 35828 129802 36148 145796
rect 65888 156044 66208 156860
rect 65888 155988 65916 156044
rect 65972 155988 66020 156044
rect 66076 155988 66124 156044
rect 66180 155988 66208 156044
rect 65888 154476 66208 155988
rect 65888 154420 65916 154476
rect 65972 154420 66020 154476
rect 66076 154420 66124 154476
rect 66180 154420 66208 154476
rect 65888 152908 66208 154420
rect 65888 152852 65916 152908
rect 65972 152852 66020 152908
rect 66076 152852 66124 152908
rect 66180 152852 66208 152908
rect 65888 151340 66208 152852
rect 65888 151284 65916 151340
rect 65972 151284 66020 151340
rect 66076 151284 66124 151340
rect 66180 151284 66208 151340
rect 65888 149772 66208 151284
rect 65888 149716 65916 149772
rect 65972 149716 66020 149772
rect 66076 149716 66124 149772
rect 66180 149716 66208 149772
rect 65888 148204 66208 149716
rect 65888 148148 65916 148204
rect 65972 148148 66020 148204
rect 66076 148148 66124 148204
rect 66180 148148 66208 148204
rect 65888 146636 66208 148148
rect 65888 146580 65916 146636
rect 65972 146580 66020 146636
rect 66076 146580 66124 146636
rect 66180 146580 66208 146636
rect 65888 145068 66208 146580
rect 65888 145012 65916 145068
rect 65972 145012 66020 145068
rect 66076 145012 66124 145068
rect 66180 145012 66208 145068
rect 65888 142955 66208 145012
rect 66548 156828 66868 156860
rect 66548 156772 66576 156828
rect 66632 156772 66680 156828
rect 66736 156772 66784 156828
rect 66840 156772 66868 156828
rect 66548 155260 66868 156772
rect 66548 155204 66576 155260
rect 66632 155204 66680 155260
rect 66736 155204 66784 155260
rect 66840 155204 66868 155260
rect 66548 153692 66868 155204
rect 66548 153636 66576 153692
rect 66632 153636 66680 153692
rect 66736 153636 66784 153692
rect 66840 153636 66868 153692
rect 66548 152124 66868 153636
rect 66548 152068 66576 152124
rect 66632 152068 66680 152124
rect 66736 152068 66784 152124
rect 66840 152068 66868 152124
rect 66548 150556 66868 152068
rect 66548 150500 66576 150556
rect 66632 150500 66680 150556
rect 66736 150500 66784 150556
rect 66840 150500 66868 150556
rect 66548 148988 66868 150500
rect 66548 148932 66576 148988
rect 66632 148932 66680 148988
rect 66736 148932 66784 148988
rect 66840 148932 66868 148988
rect 66548 147420 66868 148932
rect 66548 147364 66576 147420
rect 66632 147364 66680 147420
rect 66736 147364 66784 147420
rect 66840 147364 66868 147420
rect 66548 145852 66868 147364
rect 66548 145796 66576 145852
rect 66632 145796 66680 145852
rect 66736 145796 66784 145852
rect 66840 145796 66868 145852
rect 35828 129746 35856 129802
rect 35912 129746 35960 129802
rect 36016 129746 36064 129802
rect 36120 129746 36148 129802
rect 35828 129698 36148 129746
rect 35828 129642 35856 129698
rect 35912 129642 35960 129698
rect 36016 129642 36064 129698
rect 36120 129642 36148 129698
rect 35828 129594 36148 129642
rect 35828 129538 35856 129594
rect 35912 129538 35960 129594
rect 36016 129538 36064 129594
rect 36120 129538 36148 129594
rect 35828 99166 36148 129538
rect 48518 129802 48594 129830
rect 48518 129746 48528 129802
rect 48584 129746 48594 129802
rect 48518 129698 48594 129746
rect 48518 129642 48528 129698
rect 48584 129642 48594 129698
rect 48518 129594 48594 129642
rect 48518 129538 48528 129594
rect 48584 129538 48594 129594
rect 48518 129510 48594 129538
rect 49952 129802 50028 129830
rect 49952 129746 49962 129802
rect 50018 129746 50028 129802
rect 49952 129698 50028 129746
rect 49952 129642 49962 129698
rect 50018 129642 50028 129698
rect 49952 129594 50028 129642
rect 49952 129538 49962 129594
rect 50018 129538 50028 129594
rect 49952 129510 50028 129538
rect 51404 129802 51480 129830
rect 51404 129746 51414 129802
rect 51470 129746 51480 129802
rect 51404 129698 51480 129746
rect 51404 129642 51414 129698
rect 51470 129642 51480 129698
rect 51404 129594 51480 129642
rect 51404 129538 51414 129594
rect 51470 129538 51480 129594
rect 51404 129510 51480 129538
rect 54656 129802 54732 129830
rect 54656 129746 54666 129802
rect 54722 129746 54732 129802
rect 54656 129698 54732 129746
rect 54656 129642 54666 129698
rect 54722 129642 54732 129698
rect 54656 129594 54732 129642
rect 54656 129538 54666 129594
rect 54722 129538 54732 129594
rect 54656 129510 54732 129538
rect 65722 129802 65798 129830
rect 65722 129746 65732 129802
rect 65788 129746 65798 129802
rect 65722 129698 65798 129746
rect 65722 129642 65732 129698
rect 65788 129642 65798 129698
rect 65722 129594 65798 129642
rect 65722 129538 65732 129594
rect 65788 129538 65798 129594
rect 65722 129510 65798 129538
rect 66548 129802 66868 145796
rect 66548 129746 66576 129802
rect 66632 129746 66680 129802
rect 66736 129746 66784 129802
rect 66840 129746 66868 129802
rect 66548 129698 66868 129746
rect 66548 129642 66576 129698
rect 66632 129642 66680 129698
rect 66736 129642 66784 129698
rect 66840 129642 66868 129698
rect 66548 129594 66868 129642
rect 66548 129538 66576 129594
rect 66632 129538 66680 129594
rect 66736 129538 66784 129594
rect 66840 129538 66868 129594
rect 49588 129142 49664 129170
rect 49588 129086 49598 129142
rect 49654 129086 49664 129142
rect 49588 129038 49664 129086
rect 49588 128982 49598 129038
rect 49654 128982 49664 129038
rect 49588 128934 49664 128982
rect 49588 128878 49598 128934
rect 49654 128878 49664 128934
rect 49588 128850 49664 128878
rect 50588 129142 50664 129170
rect 50588 129086 50598 129142
rect 50654 129086 50664 129142
rect 50588 129038 50664 129086
rect 50588 128982 50598 129038
rect 50654 128982 50664 129038
rect 50588 128934 50664 128982
rect 50588 128878 50598 128934
rect 50654 128878 50664 128934
rect 50588 128850 50664 128878
rect 52029 129142 52105 129170
rect 52029 129086 52039 129142
rect 52095 129086 52105 129142
rect 52029 129038 52105 129086
rect 52029 128982 52039 129038
rect 52095 128982 52105 129038
rect 52029 128934 52105 128982
rect 52029 128878 52039 128934
rect 52095 128878 52105 128934
rect 52029 128850 52105 128878
rect 60816 129142 60892 129170
rect 60816 129086 60826 129142
rect 60882 129086 60892 129142
rect 60816 129038 60892 129086
rect 60816 128982 60826 129038
rect 60882 128982 60892 129038
rect 60816 128934 60892 128982
rect 60816 128878 60826 128934
rect 60882 128878 60892 128934
rect 60816 128850 60892 128878
rect 65286 129142 65362 129170
rect 65286 129086 65296 129142
rect 65352 129086 65362 129142
rect 65286 129038 65362 129086
rect 65286 128982 65296 129038
rect 65352 128982 65362 129038
rect 65286 128934 65362 128982
rect 65286 128878 65296 128934
rect 65352 128878 65362 128934
rect 65286 128850 65362 128878
rect 35828 99110 35856 99166
rect 35912 99110 35960 99166
rect 36016 99110 36064 99166
rect 36120 99110 36148 99166
rect 35828 99062 36148 99110
rect 35828 99006 35856 99062
rect 35912 99006 35960 99062
rect 36016 99006 36064 99062
rect 36120 99006 36148 99062
rect 35828 98958 36148 99006
rect 35828 98902 35856 98958
rect 35912 98902 35960 98958
rect 36016 98902 36064 98958
rect 36120 98902 36148 98958
rect 35828 68530 36148 98902
rect 48518 99166 48594 99194
rect 48518 99110 48528 99166
rect 48584 99110 48594 99166
rect 48518 99062 48594 99110
rect 48518 99006 48528 99062
rect 48584 99006 48594 99062
rect 48518 98958 48594 99006
rect 48518 98902 48528 98958
rect 48584 98902 48594 98958
rect 48518 98874 48594 98902
rect 49952 99166 50028 99194
rect 49952 99110 49962 99166
rect 50018 99110 50028 99166
rect 49952 99062 50028 99110
rect 49952 99006 49962 99062
rect 50018 99006 50028 99062
rect 49952 98958 50028 99006
rect 49952 98902 49962 98958
rect 50018 98902 50028 98958
rect 49952 98874 50028 98902
rect 51404 99166 51480 99194
rect 51404 99110 51414 99166
rect 51470 99110 51480 99166
rect 51404 99062 51480 99110
rect 51404 99006 51414 99062
rect 51470 99006 51480 99062
rect 51404 98958 51480 99006
rect 51404 98902 51414 98958
rect 51470 98902 51480 98958
rect 51404 98874 51480 98902
rect 54656 99166 54732 99194
rect 54656 99110 54666 99166
rect 54722 99110 54732 99166
rect 54656 99062 54732 99110
rect 54656 99006 54666 99062
rect 54722 99006 54732 99062
rect 54656 98958 54732 99006
rect 54656 98902 54666 98958
rect 54722 98902 54732 98958
rect 54656 98874 54732 98902
rect 65722 99166 65798 99194
rect 65722 99110 65732 99166
rect 65788 99110 65798 99166
rect 65722 99062 65798 99110
rect 65722 99006 65732 99062
rect 65788 99006 65798 99062
rect 65722 98958 65798 99006
rect 65722 98902 65732 98958
rect 65788 98902 65798 98958
rect 65722 98874 65798 98902
rect 66548 99166 66868 129538
rect 66548 99110 66576 99166
rect 66632 99110 66680 99166
rect 66736 99110 66784 99166
rect 66840 99110 66868 99166
rect 66548 99062 66868 99110
rect 66548 99006 66576 99062
rect 66632 99006 66680 99062
rect 66736 99006 66784 99062
rect 66840 99006 66868 99062
rect 66548 98958 66868 99006
rect 66548 98902 66576 98958
rect 66632 98902 66680 98958
rect 66736 98902 66784 98958
rect 66840 98902 66868 98958
rect 49588 98506 49664 98534
rect 49588 98450 49598 98506
rect 49654 98450 49664 98506
rect 49588 98402 49664 98450
rect 49588 98346 49598 98402
rect 49654 98346 49664 98402
rect 49588 98298 49664 98346
rect 49588 98242 49598 98298
rect 49654 98242 49664 98298
rect 49588 98214 49664 98242
rect 50588 98506 50664 98534
rect 50588 98450 50598 98506
rect 50654 98450 50664 98506
rect 50588 98402 50664 98450
rect 50588 98346 50598 98402
rect 50654 98346 50664 98402
rect 50588 98298 50664 98346
rect 50588 98242 50598 98298
rect 50654 98242 50664 98298
rect 50588 98214 50664 98242
rect 52029 98506 52105 98534
rect 52029 98450 52039 98506
rect 52095 98450 52105 98506
rect 52029 98402 52105 98450
rect 52029 98346 52039 98402
rect 52095 98346 52105 98402
rect 52029 98298 52105 98346
rect 52029 98242 52039 98298
rect 52095 98242 52105 98298
rect 52029 98214 52105 98242
rect 60816 98506 60892 98534
rect 60816 98450 60826 98506
rect 60882 98450 60892 98506
rect 60816 98402 60892 98450
rect 60816 98346 60826 98402
rect 60882 98346 60892 98402
rect 60816 98298 60892 98346
rect 60816 98242 60826 98298
rect 60882 98242 60892 98298
rect 60816 98214 60892 98242
rect 65286 98506 65362 98534
rect 65286 98450 65296 98506
rect 65352 98450 65362 98506
rect 65286 98402 65362 98450
rect 65286 98346 65296 98402
rect 65352 98346 65362 98402
rect 65286 98298 65362 98346
rect 65286 98242 65296 98298
rect 65352 98242 65362 98298
rect 65286 98214 65362 98242
rect 35828 68474 35856 68530
rect 35912 68474 35960 68530
rect 36016 68474 36064 68530
rect 36120 68474 36148 68530
rect 48518 68530 48594 68558
rect 35828 68426 36148 68474
rect 35828 68370 35856 68426
rect 35912 68370 35960 68426
rect 36016 68370 36064 68426
rect 36120 68370 36148 68426
rect 44552 68459 44628 68520
rect 44552 68403 44562 68459
rect 44618 68403 44628 68459
rect 35828 68322 36148 68370
rect 35828 68266 35856 68322
rect 35912 68266 35960 68322
rect 36016 68266 36064 68322
rect 36120 68266 36148 68322
rect 35828 37894 36148 68266
rect 42572 68341 42648 68388
rect 42572 68285 42582 68341
rect 42638 68285 42648 68341
rect 42572 68238 42648 68285
rect 44552 68355 44628 68403
rect 44552 68299 44562 68355
rect 44618 68299 44628 68355
rect 44552 68238 44628 68299
rect 48518 68474 48528 68530
rect 48584 68474 48594 68530
rect 48518 68426 48594 68474
rect 48518 68370 48528 68426
rect 48584 68370 48594 68426
rect 48518 68322 48594 68370
rect 48518 68266 48528 68322
rect 48584 68266 48594 68322
rect 48518 68238 48594 68266
rect 49952 68530 50028 68558
rect 49952 68474 49962 68530
rect 50018 68474 50028 68530
rect 49952 68426 50028 68474
rect 49952 68370 49962 68426
rect 50018 68370 50028 68426
rect 49952 68322 50028 68370
rect 49952 68266 49962 68322
rect 50018 68266 50028 68322
rect 49952 68238 50028 68266
rect 51404 68530 51480 68558
rect 51404 68474 51414 68530
rect 51470 68474 51480 68530
rect 51404 68426 51480 68474
rect 51404 68370 51414 68426
rect 51470 68370 51480 68426
rect 51404 68322 51480 68370
rect 51404 68266 51414 68322
rect 51470 68266 51480 68322
rect 51404 68238 51480 68266
rect 54656 68530 54732 68558
rect 54656 68474 54666 68530
rect 54722 68474 54732 68530
rect 54656 68426 54732 68474
rect 54656 68370 54666 68426
rect 54722 68370 54732 68426
rect 54656 68322 54732 68370
rect 54656 68266 54666 68322
rect 54722 68266 54732 68322
rect 54656 68238 54732 68266
rect 65722 68530 65798 68558
rect 65722 68474 65732 68530
rect 65788 68474 65798 68530
rect 65722 68426 65798 68474
rect 65722 68370 65732 68426
rect 65788 68370 65798 68426
rect 65722 68322 65798 68370
rect 65722 68266 65732 68322
rect 65788 68266 65798 68322
rect 65722 68238 65798 68266
rect 66548 68530 66868 98902
rect 66548 68474 66576 68530
rect 66632 68474 66680 68530
rect 66736 68474 66784 68530
rect 66840 68474 66868 68530
rect 66548 68426 66868 68474
rect 66548 68370 66576 68426
rect 66632 68370 66680 68426
rect 66736 68370 66784 68426
rect 66840 68370 66868 68426
rect 66548 68322 66868 68370
rect 66548 68266 66576 68322
rect 66632 68266 66680 68322
rect 66736 68266 66784 68322
rect 66840 68266 66868 68322
rect 44684 67855 44760 67898
rect 44684 67799 44694 67855
rect 44750 67799 44760 67855
rect 44684 67751 44760 67799
rect 44684 67695 44694 67751
rect 44750 67695 44760 67751
rect 44684 67652 44760 67695
rect 46004 67855 46080 67898
rect 46004 67799 46014 67855
rect 46070 67799 46080 67855
rect 46004 67751 46080 67799
rect 46004 67695 46014 67751
rect 46070 67695 46080 67751
rect 46004 67652 46080 67695
rect 49588 67870 49664 67898
rect 49588 67814 49598 67870
rect 49654 67814 49664 67870
rect 49588 67766 49664 67814
rect 49588 67710 49598 67766
rect 49654 67710 49664 67766
rect 49588 67662 49664 67710
rect 49588 67606 49598 67662
rect 49654 67606 49664 67662
rect 49588 67578 49664 67606
rect 50588 67870 50664 67898
rect 50588 67814 50598 67870
rect 50654 67814 50664 67870
rect 50588 67766 50664 67814
rect 50588 67710 50598 67766
rect 50654 67710 50664 67766
rect 50588 67662 50664 67710
rect 50588 67606 50598 67662
rect 50654 67606 50664 67662
rect 50588 67578 50664 67606
rect 52029 67870 52105 67898
rect 52029 67814 52039 67870
rect 52095 67814 52105 67870
rect 52029 67766 52105 67814
rect 52029 67710 52039 67766
rect 52095 67710 52105 67766
rect 52029 67662 52105 67710
rect 52029 67606 52039 67662
rect 52095 67606 52105 67662
rect 52029 67578 52105 67606
rect 60816 67870 60892 67898
rect 60816 67814 60826 67870
rect 60882 67814 60892 67870
rect 60816 67766 60892 67814
rect 60816 67710 60826 67766
rect 60882 67710 60892 67766
rect 60816 67662 60892 67710
rect 60816 67606 60826 67662
rect 60882 67606 60892 67662
rect 60816 67578 60892 67606
rect 65286 67870 65362 67898
rect 65286 67814 65296 67870
rect 65352 67814 65362 67870
rect 65286 67766 65362 67814
rect 65286 67710 65296 67766
rect 65352 67710 65362 67766
rect 65286 67662 65362 67710
rect 65286 67606 65296 67662
rect 65352 67606 65362 67662
rect 65286 67578 65362 67606
rect 35828 37838 35856 37894
rect 35912 37838 35960 37894
rect 36016 37838 36064 37894
rect 36120 37838 36148 37894
rect 35828 37790 36148 37838
rect 35828 37734 35856 37790
rect 35912 37734 35960 37790
rect 36016 37734 36064 37790
rect 36120 37734 36148 37790
rect 35828 37686 36148 37734
rect 35828 37630 35856 37686
rect 35912 37630 35960 37686
rect 36016 37630 36064 37686
rect 36120 37630 36148 37686
rect 35828 17276 36148 37630
rect 43718 37894 43794 37922
rect 43718 37838 43728 37894
rect 43784 37838 43794 37894
rect 43718 37790 43794 37838
rect 43718 37734 43728 37790
rect 43784 37734 43794 37790
rect 43718 37686 43794 37734
rect 43718 37630 43728 37686
rect 43784 37630 43794 37686
rect 43718 37602 43794 37630
rect 45960 37894 46036 37922
rect 45960 37838 45970 37894
rect 46026 37838 46036 37894
rect 45960 37790 46036 37838
rect 45960 37734 45970 37790
rect 46026 37734 46036 37790
rect 45960 37686 46036 37734
rect 45960 37630 45970 37686
rect 46026 37630 46036 37686
rect 45960 37602 46036 37630
rect 47642 37894 47718 37922
rect 47642 37838 47652 37894
rect 47708 37838 47718 37894
rect 47642 37790 47718 37838
rect 47642 37734 47652 37790
rect 47708 37734 47718 37790
rect 47642 37686 47718 37734
rect 47642 37630 47652 37686
rect 47708 37630 47718 37686
rect 47642 37602 47718 37630
rect 66548 37894 66868 68266
rect 96608 156044 96928 156860
rect 96608 155988 96636 156044
rect 96692 155988 96740 156044
rect 96796 155988 96844 156044
rect 96900 155988 96928 156044
rect 96608 154476 96928 155988
rect 96608 154420 96636 154476
rect 96692 154420 96740 154476
rect 96796 154420 96844 154476
rect 96900 154420 96928 154476
rect 96608 152908 96928 154420
rect 96608 152852 96636 152908
rect 96692 152852 96740 152908
rect 96796 152852 96844 152908
rect 96900 152852 96928 152908
rect 96608 151340 96928 152852
rect 96608 151284 96636 151340
rect 96692 151284 96740 151340
rect 96796 151284 96844 151340
rect 96900 151284 96928 151340
rect 96608 149772 96928 151284
rect 96608 149716 96636 149772
rect 96692 149716 96740 149772
rect 96796 149716 96844 149772
rect 96900 149716 96928 149772
rect 96608 148204 96928 149716
rect 96608 148148 96636 148204
rect 96692 148148 96740 148204
rect 96796 148148 96844 148204
rect 96900 148148 96928 148204
rect 96608 146636 96928 148148
rect 96608 146580 96636 146636
rect 96692 146580 96740 146636
rect 96796 146580 96844 146636
rect 96900 146580 96928 146636
rect 96608 145068 96928 146580
rect 96608 145012 96636 145068
rect 96692 145012 96740 145068
rect 96796 145012 96844 145068
rect 96900 145012 96928 145068
rect 96608 129142 96928 145012
rect 96608 129086 96636 129142
rect 96692 129086 96740 129142
rect 96796 129086 96844 129142
rect 96900 129086 96928 129142
rect 96608 129038 96928 129086
rect 96608 128982 96636 129038
rect 96692 128982 96740 129038
rect 96796 128982 96844 129038
rect 96900 128982 96928 129038
rect 96608 128934 96928 128982
rect 96608 128878 96636 128934
rect 96692 128878 96740 128934
rect 96796 128878 96844 128934
rect 96900 128878 96928 128934
rect 96608 98506 96928 128878
rect 96608 98450 96636 98506
rect 96692 98450 96740 98506
rect 96796 98450 96844 98506
rect 96900 98450 96928 98506
rect 96608 98402 96928 98450
rect 96608 98346 96636 98402
rect 96692 98346 96740 98402
rect 96796 98346 96844 98402
rect 96900 98346 96928 98402
rect 96608 98298 96928 98346
rect 96608 98242 96636 98298
rect 96692 98242 96740 98298
rect 96796 98242 96844 98298
rect 96900 98242 96928 98298
rect 96608 67870 96928 98242
rect 96608 67814 96636 67870
rect 96692 67814 96740 67870
rect 96796 67814 96844 67870
rect 96900 67814 96928 67870
rect 96608 67766 96928 67814
rect 96608 67710 96636 67766
rect 96692 67710 96740 67766
rect 96796 67710 96844 67766
rect 96900 67710 96928 67766
rect 96608 67662 96928 67710
rect 96608 67606 96636 67662
rect 96692 67606 96740 67662
rect 96796 67606 96844 67662
rect 96900 67606 96928 67662
rect 96608 39876 96928 67606
rect 97268 156828 97588 156860
rect 97268 156772 97296 156828
rect 97352 156772 97400 156828
rect 97456 156772 97504 156828
rect 97560 156772 97588 156828
rect 97268 155260 97588 156772
rect 97268 155204 97296 155260
rect 97352 155204 97400 155260
rect 97456 155204 97504 155260
rect 97560 155204 97588 155260
rect 97268 153692 97588 155204
rect 97268 153636 97296 153692
rect 97352 153636 97400 153692
rect 97456 153636 97504 153692
rect 97560 153636 97588 153692
rect 97268 152124 97588 153636
rect 97268 152068 97296 152124
rect 97352 152068 97400 152124
rect 97456 152068 97504 152124
rect 97560 152068 97588 152124
rect 97268 150556 97588 152068
rect 97268 150500 97296 150556
rect 97352 150500 97400 150556
rect 97456 150500 97504 150556
rect 97560 150500 97588 150556
rect 97268 148988 97588 150500
rect 97268 148932 97296 148988
rect 97352 148932 97400 148988
rect 97456 148932 97504 148988
rect 97560 148932 97588 148988
rect 97268 147420 97588 148932
rect 97268 147364 97296 147420
rect 97352 147364 97400 147420
rect 97456 147364 97504 147420
rect 97560 147364 97588 147420
rect 97268 145852 97588 147364
rect 97268 145796 97296 145852
rect 97352 145796 97400 145852
rect 97456 145796 97504 145852
rect 97560 145796 97588 145852
rect 97268 129802 97588 145796
rect 97268 129746 97296 129802
rect 97352 129746 97400 129802
rect 97456 129746 97504 129802
rect 97560 129746 97588 129802
rect 97268 129698 97588 129746
rect 97268 129642 97296 129698
rect 97352 129642 97400 129698
rect 97456 129642 97504 129698
rect 97560 129642 97588 129698
rect 97268 129594 97588 129642
rect 97268 129538 97296 129594
rect 97352 129538 97400 129594
rect 97456 129538 97504 129594
rect 97560 129538 97588 129594
rect 97268 99166 97588 129538
rect 97268 99110 97296 99166
rect 97352 99110 97400 99166
rect 97456 99110 97504 99166
rect 97560 99110 97588 99166
rect 97268 99062 97588 99110
rect 97268 99006 97296 99062
rect 97352 99006 97400 99062
rect 97456 99006 97504 99062
rect 97560 99006 97588 99062
rect 97268 98958 97588 99006
rect 97268 98902 97296 98958
rect 97352 98902 97400 98958
rect 97456 98902 97504 98958
rect 97560 98902 97588 98958
rect 97268 68530 97588 98902
rect 97268 68474 97296 68530
rect 97352 68474 97400 68530
rect 97456 68474 97504 68530
rect 97560 68474 97588 68530
rect 97268 68426 97588 68474
rect 97268 68370 97296 68426
rect 97352 68370 97400 68426
rect 97456 68370 97504 68426
rect 97560 68370 97588 68426
rect 97268 68322 97588 68370
rect 97268 68266 97296 68322
rect 97352 68266 97400 68322
rect 97456 68266 97504 68322
rect 97560 68266 97588 68322
rect 66548 37838 66576 37894
rect 66632 37838 66680 37894
rect 66736 37838 66784 37894
rect 66840 37838 66868 37894
rect 66548 37790 66868 37838
rect 66548 37734 66576 37790
rect 66632 37734 66680 37790
rect 66736 37734 66784 37790
rect 66840 37734 66868 37790
rect 66548 37686 66868 37734
rect 66548 37630 66576 37686
rect 66632 37630 66680 37686
rect 66736 37630 66784 37686
rect 66840 37630 66868 37686
rect 40064 37234 40140 37262
rect 40064 37178 40074 37234
rect 40130 37178 40140 37234
rect 40064 37130 40140 37178
rect 40064 37074 40074 37130
rect 40130 37074 40140 37130
rect 40064 37026 40140 37074
rect 40064 36970 40074 37026
rect 40130 36970 40140 37026
rect 40064 36942 40140 36970
rect 44374 37234 44450 37262
rect 44374 37178 44384 37234
rect 44440 37178 44450 37234
rect 44374 37130 44450 37178
rect 44374 37074 44384 37130
rect 44440 37074 44450 37130
rect 44374 37026 44450 37074
rect 44374 36970 44384 37026
rect 44440 36970 44450 37026
rect 44374 36942 44450 36970
rect 47284 37234 47360 37262
rect 47284 37178 47294 37234
rect 47350 37178 47360 37234
rect 47284 37130 47360 37178
rect 47284 37074 47294 37130
rect 47350 37074 47360 37130
rect 47284 37026 47360 37074
rect 47284 36970 47294 37026
rect 47350 36970 47360 37026
rect 47284 36942 47360 36970
rect 48298 37234 48374 37262
rect 48298 37178 48308 37234
rect 48364 37178 48374 37234
rect 48298 37130 48374 37178
rect 48298 37074 48308 37130
rect 48364 37074 48374 37130
rect 48298 37026 48374 37074
rect 48298 36970 48308 37026
rect 48364 36970 48374 37026
rect 48298 36942 48374 36970
rect 66548 35384 66868 37630
rect 97268 37894 97588 68266
rect 97268 37838 97296 37894
rect 97352 37838 97400 37894
rect 97456 37838 97504 37894
rect 97560 37838 97588 37894
rect 97268 37790 97588 37838
rect 97268 37734 97296 37790
rect 97352 37734 97400 37790
rect 97456 37734 97504 37790
rect 97560 37734 97588 37790
rect 97268 37686 97588 37734
rect 97268 37630 97296 37686
rect 97352 37630 97400 37686
rect 97456 37630 97504 37686
rect 97560 37630 97588 37686
rect 97268 35384 97588 37630
rect 127328 156044 127648 156860
rect 127328 155988 127356 156044
rect 127412 155988 127460 156044
rect 127516 155988 127564 156044
rect 127620 155988 127648 156044
rect 127328 154476 127648 155988
rect 127328 154420 127356 154476
rect 127412 154420 127460 154476
rect 127516 154420 127564 154476
rect 127620 154420 127648 154476
rect 127328 152908 127648 154420
rect 127328 152852 127356 152908
rect 127412 152852 127460 152908
rect 127516 152852 127564 152908
rect 127620 152852 127648 152908
rect 127328 151340 127648 152852
rect 127328 151284 127356 151340
rect 127412 151284 127460 151340
rect 127516 151284 127564 151340
rect 127620 151284 127648 151340
rect 127328 149772 127648 151284
rect 127328 149716 127356 149772
rect 127412 149716 127460 149772
rect 127516 149716 127564 149772
rect 127620 149716 127648 149772
rect 127328 148204 127648 149716
rect 127328 148148 127356 148204
rect 127412 148148 127460 148204
rect 127516 148148 127564 148204
rect 127620 148148 127648 148204
rect 127328 146636 127648 148148
rect 127328 146580 127356 146636
rect 127412 146580 127460 146636
rect 127516 146580 127564 146636
rect 127620 146580 127648 146636
rect 127328 145068 127648 146580
rect 127328 145012 127356 145068
rect 127412 145012 127460 145068
rect 127516 145012 127564 145068
rect 127620 145012 127648 145068
rect 127328 129142 127648 145012
rect 127328 129086 127356 129142
rect 127412 129086 127460 129142
rect 127516 129086 127564 129142
rect 127620 129086 127648 129142
rect 127328 129038 127648 129086
rect 127328 128982 127356 129038
rect 127412 128982 127460 129038
rect 127516 128982 127564 129038
rect 127620 128982 127648 129038
rect 127328 128934 127648 128982
rect 127328 128878 127356 128934
rect 127412 128878 127460 128934
rect 127516 128878 127564 128934
rect 127620 128878 127648 128934
rect 127328 98506 127648 128878
rect 127328 98450 127356 98506
rect 127412 98450 127460 98506
rect 127516 98450 127564 98506
rect 127620 98450 127648 98506
rect 127328 98402 127648 98450
rect 127328 98346 127356 98402
rect 127412 98346 127460 98402
rect 127516 98346 127564 98402
rect 127620 98346 127648 98402
rect 127328 98298 127648 98346
rect 127328 98242 127356 98298
rect 127412 98242 127460 98298
rect 127516 98242 127564 98298
rect 127620 98242 127648 98298
rect 127328 67870 127648 98242
rect 127328 67814 127356 67870
rect 127412 67814 127460 67870
rect 127516 67814 127564 67870
rect 127620 67814 127648 67870
rect 127328 67766 127648 67814
rect 127328 67710 127356 67766
rect 127412 67710 127460 67766
rect 127516 67710 127564 67766
rect 127620 67710 127648 67766
rect 127328 67662 127648 67710
rect 127328 67606 127356 67662
rect 127412 67606 127460 67662
rect 127516 67606 127564 67662
rect 127620 67606 127648 67662
rect 127328 37234 127648 67606
rect 127328 37178 127356 37234
rect 127412 37178 127460 37234
rect 127516 37178 127564 37234
rect 127620 37178 127648 37234
rect 127328 37130 127648 37178
rect 127328 37074 127356 37130
rect 127412 37074 127460 37130
rect 127516 37074 127564 37130
rect 127620 37074 127648 37130
rect 127328 37026 127648 37074
rect 127328 36970 127356 37026
rect 127412 36970 127460 37026
rect 127516 36970 127564 37026
rect 127620 36970 127648 37026
rect 127328 35384 127648 36970
rect 127988 156828 128308 156860
rect 127988 156772 128016 156828
rect 128072 156772 128120 156828
rect 128176 156772 128224 156828
rect 128280 156772 128308 156828
rect 127988 155260 128308 156772
rect 127988 155204 128016 155260
rect 128072 155204 128120 155260
rect 128176 155204 128224 155260
rect 128280 155204 128308 155260
rect 127988 153692 128308 155204
rect 127988 153636 128016 153692
rect 128072 153636 128120 153692
rect 128176 153636 128224 153692
rect 128280 153636 128308 153692
rect 127988 152124 128308 153636
rect 127988 152068 128016 152124
rect 128072 152068 128120 152124
rect 128176 152068 128224 152124
rect 128280 152068 128308 152124
rect 127988 150556 128308 152068
rect 127988 150500 128016 150556
rect 128072 150500 128120 150556
rect 128176 150500 128224 150556
rect 128280 150500 128308 150556
rect 127988 148988 128308 150500
rect 127988 148932 128016 148988
rect 128072 148932 128120 148988
rect 128176 148932 128224 148988
rect 128280 148932 128308 148988
rect 127988 147420 128308 148932
rect 127988 147364 128016 147420
rect 128072 147364 128120 147420
rect 128176 147364 128224 147420
rect 128280 147364 128308 147420
rect 127988 145852 128308 147364
rect 127988 145796 128016 145852
rect 128072 145796 128120 145852
rect 128176 145796 128224 145852
rect 128280 145796 128308 145852
rect 127988 129802 128308 145796
rect 127988 129746 128016 129802
rect 128072 129746 128120 129802
rect 128176 129746 128224 129802
rect 128280 129746 128308 129802
rect 127988 129698 128308 129746
rect 127988 129642 128016 129698
rect 128072 129642 128120 129698
rect 128176 129642 128224 129698
rect 128280 129642 128308 129698
rect 127988 129594 128308 129642
rect 127988 129538 128016 129594
rect 128072 129538 128120 129594
rect 128176 129538 128224 129594
rect 128280 129538 128308 129594
rect 127988 99166 128308 129538
rect 127988 99110 128016 99166
rect 128072 99110 128120 99166
rect 128176 99110 128224 99166
rect 128280 99110 128308 99166
rect 127988 99062 128308 99110
rect 127988 99006 128016 99062
rect 128072 99006 128120 99062
rect 128176 99006 128224 99062
rect 128280 99006 128308 99062
rect 127988 98958 128308 99006
rect 127988 98902 128016 98958
rect 128072 98902 128120 98958
rect 128176 98902 128224 98958
rect 128280 98902 128308 98958
rect 127988 68530 128308 98902
rect 127988 68474 128016 68530
rect 128072 68474 128120 68530
rect 128176 68474 128224 68530
rect 128280 68474 128308 68530
rect 127988 68426 128308 68474
rect 127988 68370 128016 68426
rect 128072 68370 128120 68426
rect 128176 68370 128224 68426
rect 128280 68370 128308 68426
rect 127988 68322 128308 68370
rect 127988 68266 128016 68322
rect 128072 68266 128120 68322
rect 128176 68266 128224 68322
rect 128280 68266 128308 68322
rect 127988 37894 128308 68266
rect 158048 156044 158368 156860
rect 158048 155988 158076 156044
rect 158132 155988 158180 156044
rect 158236 155988 158284 156044
rect 158340 155988 158368 156044
rect 158048 154476 158368 155988
rect 158048 154420 158076 154476
rect 158132 154420 158180 154476
rect 158236 154420 158284 154476
rect 158340 154420 158368 154476
rect 158048 152908 158368 154420
rect 158048 152852 158076 152908
rect 158132 152852 158180 152908
rect 158236 152852 158284 152908
rect 158340 152852 158368 152908
rect 158048 151340 158368 152852
rect 158048 151284 158076 151340
rect 158132 151284 158180 151340
rect 158236 151284 158284 151340
rect 158340 151284 158368 151340
rect 158048 149772 158368 151284
rect 158048 149716 158076 149772
rect 158132 149716 158180 149772
rect 158236 149716 158284 149772
rect 158340 149716 158368 149772
rect 158048 148204 158368 149716
rect 158048 148148 158076 148204
rect 158132 148148 158180 148204
rect 158236 148148 158284 148204
rect 158340 148148 158368 148204
rect 158048 146636 158368 148148
rect 158048 146580 158076 146636
rect 158132 146580 158180 146636
rect 158236 146580 158284 146636
rect 158340 146580 158368 146636
rect 158048 145068 158368 146580
rect 158048 145012 158076 145068
rect 158132 145012 158180 145068
rect 158236 145012 158284 145068
rect 158340 145012 158368 145068
rect 158048 129142 158368 145012
rect 158048 129086 158076 129142
rect 158132 129086 158180 129142
rect 158236 129086 158284 129142
rect 158340 129086 158368 129142
rect 158048 129038 158368 129086
rect 158048 128982 158076 129038
rect 158132 128982 158180 129038
rect 158236 128982 158284 129038
rect 158340 128982 158368 129038
rect 158048 128934 158368 128982
rect 158048 128878 158076 128934
rect 158132 128878 158180 128934
rect 158236 128878 158284 128934
rect 158340 128878 158368 128934
rect 158048 98506 158368 128878
rect 158048 98450 158076 98506
rect 158132 98450 158180 98506
rect 158236 98450 158284 98506
rect 158340 98450 158368 98506
rect 158048 98402 158368 98450
rect 158048 98346 158076 98402
rect 158132 98346 158180 98402
rect 158236 98346 158284 98402
rect 158340 98346 158368 98402
rect 158048 98298 158368 98346
rect 158048 98242 158076 98298
rect 158132 98242 158180 98298
rect 158236 98242 158284 98298
rect 158340 98242 158368 98298
rect 158048 67870 158368 98242
rect 158048 67814 158076 67870
rect 158132 67814 158180 67870
rect 158236 67814 158284 67870
rect 158340 67814 158368 67870
rect 158048 67766 158368 67814
rect 158048 67710 158076 67766
rect 158132 67710 158180 67766
rect 158236 67710 158284 67766
rect 158340 67710 158368 67766
rect 158048 67662 158368 67710
rect 158048 67606 158076 67662
rect 158132 67606 158180 67662
rect 158236 67606 158284 67662
rect 158340 67606 158368 67662
rect 132972 47012 133028 47022
rect 132972 45780 133028 46956
rect 132972 45714 133028 45724
rect 156380 47012 156436 47022
rect 156380 45780 156436 46956
rect 156380 45714 156436 45724
rect 127988 37838 128016 37894
rect 128072 37838 128120 37894
rect 128176 37838 128224 37894
rect 128280 37838 128308 37894
rect 127988 37790 128308 37838
rect 127988 37734 128016 37790
rect 128072 37734 128120 37790
rect 128176 37734 128224 37790
rect 128280 37734 128308 37790
rect 127988 37686 128308 37734
rect 127988 37630 128016 37686
rect 128072 37630 128120 37686
rect 128176 37630 128224 37686
rect 128280 37630 128308 37686
rect 82348 31892 82404 31902
rect 82348 31798 82404 31836
rect 82210 31770 82404 31798
rect 82182 31742 82404 31770
rect 77196 25396 77252 25406
rect 44156 21812 44212 21822
rect 44156 21718 44212 21756
rect 54348 21812 54404 21822
rect 54348 21718 54404 21756
rect 68348 21812 68404 21822
rect 68348 21718 68404 21756
rect 75292 21812 75348 21822
rect 75292 21718 75348 21756
rect 44156 21662 44772 21718
rect 54348 21700 55188 21718
rect 54348 21662 55132 21700
rect 44716 21252 44772 21662
rect 68348 21662 68746 21718
rect 75292 21662 75478 21718
rect 55132 21634 55188 21644
rect 44716 21186 44772 21196
rect 77196 21140 77252 25340
rect 82182 25318 82238 31742
rect 125356 26068 125412 26078
rect 125412 26012 125506 26038
rect 125356 25982 125506 26012
rect 96572 25508 96628 25518
rect 96628 25452 96730 25498
rect 96572 25442 96730 25452
rect 78652 25284 78708 25294
rect 78652 21252 78708 25228
rect 82012 25290 82238 25318
rect 110908 25396 110964 25406
rect 110908 25318 110964 25340
rect 82012 25284 82210 25290
rect 82068 25262 82210 25284
rect 110908 25262 111118 25318
rect 82012 25218 82068 25228
rect 78652 21186 78708 21196
rect 77196 21074 77252 21084
rect 48300 20468 48356 20478
rect 48154 20412 48300 20458
rect 48154 20402 48356 20412
rect 67788 20468 67844 20478
rect 82460 20468 82516 20478
rect 67844 20412 67954 20458
rect 67788 20402 67954 20412
rect 82342 20412 82460 20458
rect 82342 20402 82516 20412
rect 58318 20042 58772 20098
rect 58716 19908 58772 20042
rect 58716 19842 58772 19852
rect 35828 17220 35856 17276
rect 35912 17220 35960 17276
rect 36016 17220 36064 17276
rect 36120 17220 36148 17276
rect 35828 15708 36148 17220
rect 35828 15652 35856 15708
rect 35912 15652 35960 15708
rect 36016 15652 36064 15708
rect 36120 15652 36148 15708
rect 35828 14140 36148 15652
rect 35828 14084 35856 14140
rect 35912 14084 35960 14140
rect 36016 14084 36064 14140
rect 36120 14084 36148 14140
rect 35828 12572 36148 14084
rect 35828 12516 35856 12572
rect 35912 12516 35960 12572
rect 36016 12516 36064 12572
rect 36120 12516 36148 12572
rect 35828 11004 36148 12516
rect 35828 10948 35856 11004
rect 35912 10948 35960 11004
rect 36016 10948 36064 11004
rect 36120 10948 36148 11004
rect 35828 9436 36148 10948
rect 35828 9380 35856 9436
rect 35912 9380 35960 9436
rect 36016 9380 36064 9436
rect 36120 9380 36148 9436
rect 35828 7868 36148 9380
rect 35828 7812 35856 7868
rect 35912 7812 35960 7868
rect 36016 7812 36064 7868
rect 36120 7812 36148 7868
rect 35828 7258 36148 7812
rect 35828 7202 35856 7258
rect 35912 7202 35960 7258
rect 36016 7202 36064 7258
rect 36120 7202 36148 7258
rect 35828 7154 36148 7202
rect 35828 7098 35856 7154
rect 35912 7098 35960 7154
rect 36016 7098 36064 7154
rect 36120 7098 36148 7154
rect 35828 7050 36148 7098
rect 35828 6994 35856 7050
rect 35912 6994 35960 7050
rect 36016 6994 36064 7050
rect 36120 6994 36148 7050
rect 35828 6300 36148 6994
rect 35828 6244 35856 6300
rect 35912 6244 35960 6300
rect 36016 6244 36064 6300
rect 36120 6244 36148 6300
rect 35828 4732 36148 6244
rect 35828 4676 35856 4732
rect 35912 4676 35960 4732
rect 36016 4676 36064 4732
rect 36120 4676 36148 4732
rect 35828 3164 36148 4676
rect 35828 3108 35856 3164
rect 35912 3108 35960 3164
rect 36016 3108 36064 3164
rect 36120 3108 36148 3164
rect 35828 3076 36148 3108
rect 65888 16492 66208 20065
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 6598 66208 7028
rect 65888 6542 65916 6598
rect 65972 6542 66020 6598
rect 66076 6542 66124 6598
rect 66180 6542 66208 6598
rect 65888 6494 66208 6542
rect 65888 6438 65916 6494
rect 65972 6438 66020 6494
rect 66076 6438 66124 6494
rect 66180 6438 66208 6494
rect 65888 6390 66208 6438
rect 65888 6334 65916 6390
rect 65972 6334 66020 6390
rect 66076 6334 66124 6390
rect 66180 6334 66208 6390
rect 65888 5516 66208 6334
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 66548 17276 66868 20065
rect 66548 17220 66576 17276
rect 66632 17220 66680 17276
rect 66736 17220 66784 17276
rect 66840 17220 66868 17276
rect 66548 15708 66868 17220
rect 77308 18452 77364 18462
rect 77308 17108 77364 18396
rect 77308 17042 77364 17052
rect 78876 17108 78932 20098
rect 78876 17042 78932 17052
rect 66548 15652 66576 15708
rect 66632 15652 66680 15708
rect 66736 15652 66784 15708
rect 66840 15652 66868 15708
rect 66548 14140 66868 15652
rect 66548 14084 66576 14140
rect 66632 14084 66680 14140
rect 66736 14084 66784 14140
rect 66840 14084 66868 14140
rect 66548 12572 66868 14084
rect 66548 12516 66576 12572
rect 66632 12516 66680 12572
rect 66736 12516 66784 12572
rect 66840 12516 66868 12572
rect 66548 11004 66868 12516
rect 66548 10948 66576 11004
rect 66632 10948 66680 11004
rect 66736 10948 66784 11004
rect 66840 10948 66868 11004
rect 66548 9436 66868 10948
rect 66548 9380 66576 9436
rect 66632 9380 66680 9436
rect 66736 9380 66784 9436
rect 66840 9380 66868 9436
rect 66548 7868 66868 9380
rect 66548 7812 66576 7868
rect 66632 7812 66680 7868
rect 66736 7812 66784 7868
rect 66840 7812 66868 7868
rect 66548 7258 66868 7812
rect 66548 7202 66576 7258
rect 66632 7202 66680 7258
rect 66736 7202 66784 7258
rect 66840 7202 66868 7258
rect 66548 7154 66868 7202
rect 66548 7098 66576 7154
rect 66632 7098 66680 7154
rect 66736 7098 66784 7154
rect 66840 7098 66868 7154
rect 66548 7050 66868 7098
rect 66548 6994 66576 7050
rect 66632 6994 66680 7050
rect 66736 6994 66784 7050
rect 66840 6994 66868 7050
rect 66548 6300 66868 6994
rect 66548 6244 66576 6300
rect 66632 6244 66680 6300
rect 66736 6244 66784 6300
rect 66840 6244 66868 6300
rect 66548 4732 66868 6244
rect 66548 4676 66576 4732
rect 66632 4676 66680 4732
rect 66736 4676 66784 4732
rect 66840 4676 66868 4732
rect 66548 3164 66868 4676
rect 66548 3108 66576 3164
rect 66632 3108 66680 3164
rect 66736 3108 66784 3164
rect 66840 3108 66868 3164
rect 66548 3076 66868 3108
rect 96608 16492 96928 17888
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 6598 96928 7028
rect 96608 6542 96636 6598
rect 96692 6542 96740 6598
rect 96796 6542 96844 6598
rect 96900 6542 96928 6598
rect 96608 6494 96928 6542
rect 96608 6438 96636 6494
rect 96692 6438 96740 6494
rect 96796 6438 96844 6494
rect 96900 6438 96928 6494
rect 96608 6390 96928 6438
rect 96608 6334 96636 6390
rect 96692 6334 96740 6390
rect 96796 6334 96844 6390
rect 96900 6334 96928 6390
rect 96608 5516 96928 6334
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 97268 17276 97588 21056
rect 97268 17220 97296 17276
rect 97352 17220 97400 17276
rect 97456 17220 97504 17276
rect 97560 17220 97588 17276
rect 97268 15708 97588 17220
rect 97268 15652 97296 15708
rect 97352 15652 97400 15708
rect 97456 15652 97504 15708
rect 97560 15652 97588 15708
rect 97268 14140 97588 15652
rect 97268 14084 97296 14140
rect 97352 14084 97400 14140
rect 97456 14084 97504 14140
rect 97560 14084 97588 14140
rect 97268 12572 97588 14084
rect 97268 12516 97296 12572
rect 97352 12516 97400 12572
rect 97456 12516 97504 12572
rect 97560 12516 97588 12572
rect 97268 11004 97588 12516
rect 97268 10948 97296 11004
rect 97352 10948 97400 11004
rect 97456 10948 97504 11004
rect 97560 10948 97588 11004
rect 97268 9436 97588 10948
rect 97268 9380 97296 9436
rect 97352 9380 97400 9436
rect 97456 9380 97504 9436
rect 97560 9380 97588 9436
rect 97268 7868 97588 9380
rect 97268 7812 97296 7868
rect 97352 7812 97400 7868
rect 97456 7812 97504 7868
rect 97560 7812 97588 7868
rect 97268 7258 97588 7812
rect 97268 7202 97296 7258
rect 97352 7202 97400 7258
rect 97456 7202 97504 7258
rect 97560 7202 97588 7258
rect 97268 7154 97588 7202
rect 97268 7098 97296 7154
rect 97352 7098 97400 7154
rect 97456 7098 97504 7154
rect 97560 7098 97588 7154
rect 97268 7050 97588 7098
rect 97268 6994 97296 7050
rect 97352 6994 97400 7050
rect 97456 6994 97504 7050
rect 97560 6994 97588 7050
rect 97268 6300 97588 6994
rect 97268 6244 97296 6300
rect 97352 6244 97400 6300
rect 97456 6244 97504 6300
rect 97560 6244 97588 6300
rect 97268 4732 97588 6244
rect 97268 4676 97296 4732
rect 97352 4676 97400 4732
rect 97456 4676 97504 4732
rect 97560 4676 97588 4732
rect 97268 3164 97588 4676
rect 97268 3108 97296 3164
rect 97352 3108 97400 3164
rect 97456 3108 97504 3164
rect 97560 3108 97588 3164
rect 97268 3076 97588 3108
rect 127328 16492 127648 21188
rect 127328 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127648 16492
rect 127328 14924 127648 16436
rect 127328 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127648 14924
rect 127328 13356 127648 14868
rect 127328 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127648 13356
rect 127328 11788 127648 13300
rect 127328 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127648 11788
rect 127328 10220 127648 11732
rect 127328 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127648 10220
rect 127328 8652 127648 10164
rect 127328 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127648 8652
rect 127328 7084 127648 8596
rect 127328 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127648 7084
rect 127328 6598 127648 7028
rect 127328 6542 127356 6598
rect 127412 6542 127460 6598
rect 127516 6542 127564 6598
rect 127620 6542 127648 6598
rect 127328 6494 127648 6542
rect 127328 6438 127356 6494
rect 127412 6438 127460 6494
rect 127516 6438 127564 6494
rect 127620 6438 127648 6494
rect 127328 6390 127648 6438
rect 127328 6334 127356 6390
rect 127412 6334 127460 6390
rect 127516 6334 127564 6390
rect 127620 6334 127648 6390
rect 127328 5516 127648 6334
rect 127328 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127648 5516
rect 127328 3948 127648 5460
rect 127328 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127648 3948
rect 127328 3076 127648 3892
rect 127988 17276 128308 37630
rect 130880 37234 130956 37262
rect 130880 37178 130890 37234
rect 130946 37178 130956 37234
rect 130880 37130 130956 37178
rect 130880 37074 130890 37130
rect 130946 37074 130956 37130
rect 130880 37026 130956 37074
rect 130880 36970 130890 37026
rect 130946 36970 130956 37026
rect 130880 36942 130956 36970
rect 158048 37234 158368 67606
rect 158048 37178 158076 37234
rect 158132 37178 158180 37234
rect 158236 37178 158284 37234
rect 158340 37178 158368 37234
rect 158048 37130 158368 37178
rect 158048 37074 158076 37130
rect 158132 37074 158180 37130
rect 158236 37074 158284 37130
rect 158340 37074 158368 37130
rect 158048 37026 158368 37074
rect 158048 36970 158076 37026
rect 158132 36970 158180 37026
rect 158236 36970 158284 37026
rect 158340 36970 158368 37026
rect 154700 27860 154756 27870
rect 139894 26180 140084 26218
rect 139894 26162 140028 26180
rect 140028 26114 140084 26124
rect 154700 26180 154756 27804
rect 154700 26114 154756 26124
rect 155148 27748 155204 27758
rect 154812 26068 154868 26078
rect 154252 20468 154308 20478
rect 154150 20412 154252 20458
rect 154150 20402 154308 20412
rect 127988 17220 128016 17276
rect 128072 17220 128120 17276
rect 128176 17220 128224 17276
rect 128280 17220 128308 17276
rect 127988 15708 128308 17220
rect 154812 16884 154868 26012
rect 155148 26068 155204 27692
rect 155148 26002 155204 26012
rect 154812 16818 154868 16828
rect 127988 15652 128016 15708
rect 128072 15652 128120 15708
rect 128176 15652 128224 15708
rect 128280 15652 128308 15708
rect 127988 14140 128308 15652
rect 127988 14084 128016 14140
rect 128072 14084 128120 14140
rect 128176 14084 128224 14140
rect 128280 14084 128308 14140
rect 127988 12572 128308 14084
rect 127988 12516 128016 12572
rect 128072 12516 128120 12572
rect 128176 12516 128224 12572
rect 128280 12516 128308 12572
rect 127988 11004 128308 12516
rect 127988 10948 128016 11004
rect 128072 10948 128120 11004
rect 128176 10948 128224 11004
rect 128280 10948 128308 11004
rect 127988 9436 128308 10948
rect 127988 9380 128016 9436
rect 128072 9380 128120 9436
rect 128176 9380 128224 9436
rect 128280 9380 128308 9436
rect 127988 7868 128308 9380
rect 127988 7812 128016 7868
rect 128072 7812 128120 7868
rect 128176 7812 128224 7868
rect 128280 7812 128308 7868
rect 127988 7258 128308 7812
rect 127988 7202 128016 7258
rect 128072 7202 128120 7258
rect 128176 7202 128224 7258
rect 128280 7202 128308 7258
rect 127988 7154 128308 7202
rect 127988 7098 128016 7154
rect 128072 7098 128120 7154
rect 128176 7098 128224 7154
rect 128280 7098 128308 7154
rect 127988 7050 128308 7098
rect 127988 6994 128016 7050
rect 128072 6994 128120 7050
rect 128176 6994 128224 7050
rect 128280 6994 128308 7050
rect 127988 6300 128308 6994
rect 127988 6244 128016 6300
rect 128072 6244 128120 6300
rect 128176 6244 128224 6300
rect 128280 6244 128308 6300
rect 127988 4732 128308 6244
rect 127988 4676 128016 4732
rect 128072 4676 128120 4732
rect 128176 4676 128224 4732
rect 128280 4676 128308 4732
rect 127988 3164 128308 4676
rect 127988 3108 128016 3164
rect 128072 3108 128120 3164
rect 128176 3108 128224 3164
rect 128280 3108 128308 3164
rect 127988 3076 128308 3108
rect 158048 16492 158368 36970
rect 158048 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158368 16492
rect 158048 14924 158368 16436
rect 158048 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158368 14924
rect 158048 13356 158368 14868
rect 158048 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158368 13356
rect 158048 11788 158368 13300
rect 158048 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158368 11788
rect 158048 10220 158368 11732
rect 158048 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158368 10220
rect 158048 8652 158368 10164
rect 158048 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158368 8652
rect 158048 7084 158368 8596
rect 158048 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158368 7084
rect 158048 6598 158368 7028
rect 158048 6542 158076 6598
rect 158132 6542 158180 6598
rect 158236 6542 158284 6598
rect 158340 6542 158368 6598
rect 158048 6494 158368 6542
rect 158048 6438 158076 6494
rect 158132 6438 158180 6494
rect 158236 6438 158284 6494
rect 158340 6438 158368 6494
rect 158048 6390 158368 6438
rect 158048 6334 158076 6390
rect 158132 6334 158180 6390
rect 158236 6334 158284 6390
rect 158340 6334 158368 6390
rect 158048 5516 158368 6334
rect 158048 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158368 5516
rect 158048 3948 158368 5460
rect 158048 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158368 3948
rect 158048 3076 158368 3892
rect 158708 156828 159028 156860
rect 158708 156772 158736 156828
rect 158792 156772 158840 156828
rect 158896 156772 158944 156828
rect 159000 156772 159028 156828
rect 158708 155260 159028 156772
rect 158708 155204 158736 155260
rect 158792 155204 158840 155260
rect 158896 155204 158944 155260
rect 159000 155204 159028 155260
rect 158708 153692 159028 155204
rect 158708 153636 158736 153692
rect 158792 153636 158840 153692
rect 158896 153636 158944 153692
rect 159000 153636 159028 153692
rect 158708 152124 159028 153636
rect 158708 152068 158736 152124
rect 158792 152068 158840 152124
rect 158896 152068 158944 152124
rect 159000 152068 159028 152124
rect 158708 150556 159028 152068
rect 158708 150500 158736 150556
rect 158792 150500 158840 150556
rect 158896 150500 158944 150556
rect 159000 150500 159028 150556
rect 158708 148988 159028 150500
rect 158708 148932 158736 148988
rect 158792 148932 158840 148988
rect 158896 148932 158944 148988
rect 159000 148932 159028 148988
rect 158708 147420 159028 148932
rect 158708 147364 158736 147420
rect 158792 147364 158840 147420
rect 158896 147364 158944 147420
rect 159000 147364 159028 147420
rect 158708 145852 159028 147364
rect 158708 145796 158736 145852
rect 158792 145796 158840 145852
rect 158896 145796 158944 145852
rect 159000 145796 159028 145852
rect 158708 129802 159028 145796
rect 188768 156044 189088 156860
rect 188768 155988 188796 156044
rect 188852 155988 188900 156044
rect 188956 155988 189004 156044
rect 189060 155988 189088 156044
rect 188768 154476 189088 155988
rect 188768 154420 188796 154476
rect 188852 154420 188900 154476
rect 188956 154420 189004 154476
rect 189060 154420 189088 154476
rect 188768 152908 189088 154420
rect 188768 152852 188796 152908
rect 188852 152852 188900 152908
rect 188956 152852 189004 152908
rect 189060 152852 189088 152908
rect 188768 151340 189088 152852
rect 188768 151284 188796 151340
rect 188852 151284 188900 151340
rect 188956 151284 189004 151340
rect 189060 151284 189088 151340
rect 188768 149772 189088 151284
rect 188768 149716 188796 149772
rect 188852 149716 188900 149772
rect 188956 149716 189004 149772
rect 189060 149716 189088 149772
rect 188768 148204 189088 149716
rect 188768 148148 188796 148204
rect 188852 148148 188900 148204
rect 188956 148148 189004 148204
rect 189060 148148 189088 148204
rect 188768 146636 189088 148148
rect 188768 146580 188796 146636
rect 188852 146580 188900 146636
rect 188956 146580 189004 146636
rect 189060 146580 189088 146636
rect 188768 145068 189088 146580
rect 188768 145012 188796 145068
rect 188852 145012 188900 145068
rect 188956 145012 189004 145068
rect 189060 145012 189088 145068
rect 188768 143500 189088 145012
rect 188768 143444 188796 143500
rect 188852 143444 188900 143500
rect 188956 143444 189004 143500
rect 189060 143444 189088 143500
rect 188768 141932 189088 143444
rect 188768 141876 188796 141932
rect 188852 141876 188900 141932
rect 188956 141876 189004 141932
rect 189060 141876 189088 141932
rect 188768 140364 189088 141876
rect 188768 140308 188796 140364
rect 188852 140308 188900 140364
rect 188956 140308 189004 140364
rect 189060 140308 189088 140364
rect 188768 138796 189088 140308
rect 188768 138740 188796 138796
rect 188852 138740 188900 138796
rect 188956 138740 189004 138796
rect 189060 138740 189088 138796
rect 188768 137228 189088 138740
rect 188768 137172 188796 137228
rect 188852 137172 188900 137228
rect 188956 137172 189004 137228
rect 189060 137172 189088 137228
rect 188768 135660 189088 137172
rect 188768 135604 188796 135660
rect 188852 135604 188900 135660
rect 188956 135604 189004 135660
rect 189060 135604 189088 135660
rect 188768 134092 189088 135604
rect 188768 134036 188796 134092
rect 188852 134036 188900 134092
rect 188956 134036 189004 134092
rect 189060 134036 189088 134092
rect 188768 132524 189088 134036
rect 188768 132468 188796 132524
rect 188852 132468 188900 132524
rect 188956 132468 189004 132524
rect 189060 132468 189088 132524
rect 188768 130956 189088 132468
rect 188768 130900 188796 130956
rect 188852 130900 188900 130956
rect 188956 130900 189004 130956
rect 189060 130900 189088 130956
rect 158708 129746 158736 129802
rect 158792 129746 158840 129802
rect 158896 129746 158944 129802
rect 159000 129746 159028 129802
rect 158708 129698 159028 129746
rect 158708 129642 158736 129698
rect 158792 129642 158840 129698
rect 158896 129642 158944 129698
rect 159000 129642 159028 129698
rect 158708 129594 159028 129642
rect 158708 129538 158736 129594
rect 158792 129538 158840 129594
rect 158896 129538 158944 129594
rect 159000 129538 159028 129594
rect 158708 99166 159028 129538
rect 184012 129802 184088 129830
rect 184012 129746 184022 129802
rect 184078 129746 184088 129802
rect 184012 129698 184088 129746
rect 184012 129642 184022 129698
rect 184078 129642 184088 129698
rect 184012 129594 184088 129642
rect 184012 129538 184022 129594
rect 184078 129538 184088 129594
rect 184012 129510 184088 129538
rect 185924 129802 186264 129830
rect 185924 129746 185962 129802
rect 186018 129746 186066 129802
rect 186122 129746 186170 129802
rect 186226 129746 186264 129802
rect 185924 129698 186264 129746
rect 185924 129642 185962 129698
rect 186018 129642 186066 129698
rect 186122 129642 186170 129698
rect 186226 129642 186264 129698
rect 185924 129594 186264 129642
rect 185924 129538 185962 129594
rect 186018 129538 186066 129594
rect 186122 129538 186170 129594
rect 186226 129538 186264 129594
rect 185924 129510 186264 129538
rect 188768 129388 189088 130900
rect 188768 129332 188796 129388
rect 188852 129332 188900 129388
rect 188956 129332 189004 129388
rect 189060 129332 189088 129388
rect 184448 129142 184524 129170
rect 184448 129086 184458 129142
rect 184514 129086 184524 129142
rect 184448 129038 184524 129086
rect 184448 128982 184458 129038
rect 184514 128982 184524 129038
rect 184448 128934 184524 128982
rect 184448 128878 184458 128934
rect 184514 128878 184524 128934
rect 184448 128850 184524 128878
rect 185264 129142 185604 129170
rect 185264 129086 185302 129142
rect 185358 129086 185406 129142
rect 185462 129086 185510 129142
rect 185566 129086 185604 129142
rect 185264 129038 185604 129086
rect 185264 128982 185302 129038
rect 185358 128982 185406 129038
rect 185462 128982 185510 129038
rect 185566 128982 185604 129038
rect 185264 128934 185604 128982
rect 185264 128878 185302 128934
rect 185358 128878 185406 128934
rect 185462 128878 185510 128934
rect 185566 128878 185604 128934
rect 185264 128850 185604 128878
rect 188768 129142 189088 129332
rect 188768 129086 188796 129142
rect 188852 129086 188900 129142
rect 188956 129086 189004 129142
rect 189060 129086 189088 129142
rect 188768 129038 189088 129086
rect 188768 128982 188796 129038
rect 188852 128982 188900 129038
rect 188956 128982 189004 129038
rect 189060 128982 189088 129038
rect 188768 128934 189088 128982
rect 188768 128878 188796 128934
rect 188852 128878 188900 128934
rect 188956 128878 189004 128934
rect 189060 128878 189088 128934
rect 188768 127820 189088 128878
rect 188768 127764 188796 127820
rect 188852 127764 188900 127820
rect 188956 127764 189004 127820
rect 189060 127764 189088 127820
rect 188768 126252 189088 127764
rect 188768 126196 188796 126252
rect 188852 126196 188900 126252
rect 188956 126196 189004 126252
rect 189060 126196 189088 126252
rect 188768 124684 189088 126196
rect 188768 124628 188796 124684
rect 188852 124628 188900 124684
rect 188956 124628 189004 124684
rect 189060 124628 189088 124684
rect 188768 123116 189088 124628
rect 188768 123060 188796 123116
rect 188852 123060 188900 123116
rect 188956 123060 189004 123116
rect 189060 123060 189088 123116
rect 188768 121548 189088 123060
rect 188768 121492 188796 121548
rect 188852 121492 188900 121548
rect 188956 121492 189004 121548
rect 189060 121492 189088 121548
rect 188768 119980 189088 121492
rect 188768 119924 188796 119980
rect 188852 119924 188900 119980
rect 188956 119924 189004 119980
rect 189060 119924 189088 119980
rect 188768 118412 189088 119924
rect 188768 118356 188796 118412
rect 188852 118356 188900 118412
rect 188956 118356 189004 118412
rect 189060 118356 189088 118412
rect 188768 116844 189088 118356
rect 188768 116788 188796 116844
rect 188852 116788 188900 116844
rect 188956 116788 189004 116844
rect 189060 116788 189088 116844
rect 188768 115276 189088 116788
rect 188768 115220 188796 115276
rect 188852 115220 188900 115276
rect 188956 115220 189004 115276
rect 189060 115220 189088 115276
rect 188768 113708 189088 115220
rect 188768 113652 188796 113708
rect 188852 113652 188900 113708
rect 188956 113652 189004 113708
rect 189060 113652 189088 113708
rect 188768 112140 189088 113652
rect 188768 112084 188796 112140
rect 188852 112084 188900 112140
rect 188956 112084 189004 112140
rect 189060 112084 189088 112140
rect 188768 110572 189088 112084
rect 188768 110516 188796 110572
rect 188852 110516 188900 110572
rect 188956 110516 189004 110572
rect 189060 110516 189088 110572
rect 188768 109004 189088 110516
rect 188768 108948 188796 109004
rect 188852 108948 188900 109004
rect 188956 108948 189004 109004
rect 189060 108948 189088 109004
rect 188768 107436 189088 108948
rect 188768 107380 188796 107436
rect 188852 107380 188900 107436
rect 188956 107380 189004 107436
rect 189060 107380 189088 107436
rect 188768 105868 189088 107380
rect 188768 105812 188796 105868
rect 188852 105812 188900 105868
rect 188956 105812 189004 105868
rect 189060 105812 189088 105868
rect 188768 104300 189088 105812
rect 188768 104244 188796 104300
rect 188852 104244 188900 104300
rect 188956 104244 189004 104300
rect 189060 104244 189088 104300
rect 188768 102732 189088 104244
rect 188768 102676 188796 102732
rect 188852 102676 188900 102732
rect 188956 102676 189004 102732
rect 189060 102676 189088 102732
rect 188768 101164 189088 102676
rect 188768 101108 188796 101164
rect 188852 101108 188900 101164
rect 188956 101108 189004 101164
rect 189060 101108 189088 101164
rect 188768 99596 189088 101108
rect 188768 99540 188796 99596
rect 188852 99540 188900 99596
rect 188956 99540 189004 99596
rect 189060 99540 189088 99596
rect 158708 99110 158736 99166
rect 158792 99110 158840 99166
rect 158896 99110 158944 99166
rect 159000 99110 159028 99166
rect 158708 99062 159028 99110
rect 158708 99006 158736 99062
rect 158792 99006 158840 99062
rect 158896 99006 158944 99062
rect 159000 99006 159028 99062
rect 158708 98958 159028 99006
rect 158708 98902 158736 98958
rect 158792 98902 158840 98958
rect 158896 98902 158944 98958
rect 159000 98902 159028 98958
rect 158708 68530 159028 98902
rect 184012 99166 184088 99194
rect 184012 99110 184022 99166
rect 184078 99110 184088 99166
rect 184012 99062 184088 99110
rect 184012 99006 184022 99062
rect 184078 99006 184088 99062
rect 184012 98958 184088 99006
rect 184012 98902 184022 98958
rect 184078 98902 184088 98958
rect 184012 98874 184088 98902
rect 185924 99166 186264 99194
rect 185924 99110 185962 99166
rect 186018 99110 186066 99166
rect 186122 99110 186170 99166
rect 186226 99110 186264 99166
rect 185924 99062 186264 99110
rect 185924 99006 185962 99062
rect 186018 99006 186066 99062
rect 186122 99006 186170 99062
rect 186226 99006 186264 99062
rect 185924 98958 186264 99006
rect 185924 98902 185962 98958
rect 186018 98902 186066 98958
rect 186122 98902 186170 98958
rect 186226 98902 186264 98958
rect 185924 98874 186264 98902
rect 184448 98506 184524 98534
rect 184448 98450 184458 98506
rect 184514 98450 184524 98506
rect 184448 98402 184524 98450
rect 184448 98346 184458 98402
rect 184514 98346 184524 98402
rect 184448 98298 184524 98346
rect 184448 98242 184458 98298
rect 184514 98242 184524 98298
rect 184448 98214 184524 98242
rect 185264 98506 185604 98534
rect 185264 98450 185302 98506
rect 185358 98450 185406 98506
rect 185462 98450 185510 98506
rect 185566 98450 185604 98506
rect 185264 98402 185604 98450
rect 185264 98346 185302 98402
rect 185358 98346 185406 98402
rect 185462 98346 185510 98402
rect 185566 98346 185604 98402
rect 185264 98298 185604 98346
rect 185264 98242 185302 98298
rect 185358 98242 185406 98298
rect 185462 98242 185510 98298
rect 185566 98242 185604 98298
rect 185264 98214 185604 98242
rect 188768 98506 189088 99540
rect 188768 98450 188796 98506
rect 188852 98450 188900 98506
rect 188956 98450 189004 98506
rect 189060 98450 189088 98506
rect 188768 98402 189088 98450
rect 188768 98346 188796 98402
rect 188852 98346 188900 98402
rect 188956 98346 189004 98402
rect 189060 98346 189088 98402
rect 188768 98298 189088 98346
rect 188768 98242 188796 98298
rect 188852 98242 188900 98298
rect 188956 98242 189004 98298
rect 189060 98242 189088 98298
rect 188768 98028 189088 98242
rect 188768 97972 188796 98028
rect 188852 97972 188900 98028
rect 188956 97972 189004 98028
rect 189060 97972 189088 98028
rect 188768 96460 189088 97972
rect 188768 96404 188796 96460
rect 188852 96404 188900 96460
rect 188956 96404 189004 96460
rect 189060 96404 189088 96460
rect 188768 94892 189088 96404
rect 188768 94836 188796 94892
rect 188852 94836 188900 94892
rect 188956 94836 189004 94892
rect 189060 94836 189088 94892
rect 188768 93324 189088 94836
rect 188768 93268 188796 93324
rect 188852 93268 188900 93324
rect 188956 93268 189004 93324
rect 189060 93268 189088 93324
rect 188768 91756 189088 93268
rect 188768 91700 188796 91756
rect 188852 91700 188900 91756
rect 188956 91700 189004 91756
rect 189060 91700 189088 91756
rect 188768 90188 189088 91700
rect 188768 90132 188796 90188
rect 188852 90132 188900 90188
rect 188956 90132 189004 90188
rect 189060 90132 189088 90188
rect 188768 88620 189088 90132
rect 188768 88564 188796 88620
rect 188852 88564 188900 88620
rect 188956 88564 189004 88620
rect 189060 88564 189088 88620
rect 188768 87052 189088 88564
rect 188768 86996 188796 87052
rect 188852 86996 188900 87052
rect 188956 86996 189004 87052
rect 189060 86996 189088 87052
rect 188768 85484 189088 86996
rect 188768 85428 188796 85484
rect 188852 85428 188900 85484
rect 188956 85428 189004 85484
rect 189060 85428 189088 85484
rect 188768 83916 189088 85428
rect 188768 83860 188796 83916
rect 188852 83860 188900 83916
rect 188956 83860 189004 83916
rect 189060 83860 189088 83916
rect 188768 82348 189088 83860
rect 188768 82292 188796 82348
rect 188852 82292 188900 82348
rect 188956 82292 189004 82348
rect 189060 82292 189088 82348
rect 188768 80780 189088 82292
rect 188768 80724 188796 80780
rect 188852 80724 188900 80780
rect 188956 80724 189004 80780
rect 189060 80724 189088 80780
rect 188768 79212 189088 80724
rect 188768 79156 188796 79212
rect 188852 79156 188900 79212
rect 188956 79156 189004 79212
rect 189060 79156 189088 79212
rect 188768 77644 189088 79156
rect 188768 77588 188796 77644
rect 188852 77588 188900 77644
rect 188956 77588 189004 77644
rect 189060 77588 189088 77644
rect 188768 76076 189088 77588
rect 188768 76020 188796 76076
rect 188852 76020 188900 76076
rect 188956 76020 189004 76076
rect 189060 76020 189088 76076
rect 188768 74508 189088 76020
rect 188768 74452 188796 74508
rect 188852 74452 188900 74508
rect 188956 74452 189004 74508
rect 189060 74452 189088 74508
rect 188768 72940 189088 74452
rect 188768 72884 188796 72940
rect 188852 72884 188900 72940
rect 188956 72884 189004 72940
rect 189060 72884 189088 72940
rect 188768 71372 189088 72884
rect 188768 71316 188796 71372
rect 188852 71316 188900 71372
rect 188956 71316 189004 71372
rect 189060 71316 189088 71372
rect 188768 69804 189088 71316
rect 188768 69748 188796 69804
rect 188852 69748 188900 69804
rect 188956 69748 189004 69804
rect 189060 69748 189088 69804
rect 158708 68474 158736 68530
rect 158792 68474 158840 68530
rect 158896 68474 158944 68530
rect 159000 68474 159028 68530
rect 158708 68426 159028 68474
rect 158708 68370 158736 68426
rect 158792 68370 158840 68426
rect 158896 68370 158944 68426
rect 159000 68370 159028 68426
rect 158708 68322 159028 68370
rect 158708 68266 158736 68322
rect 158792 68266 158840 68322
rect 158896 68266 158944 68322
rect 159000 68266 159028 68322
rect 158708 37894 159028 68266
rect 184012 68530 184088 68558
rect 184012 68474 184022 68530
rect 184078 68474 184088 68530
rect 184012 68426 184088 68474
rect 184012 68370 184022 68426
rect 184078 68370 184088 68426
rect 184012 68322 184088 68370
rect 184012 68266 184022 68322
rect 184078 68266 184088 68322
rect 184012 68238 184088 68266
rect 185924 68530 186264 68558
rect 185924 68474 185962 68530
rect 186018 68474 186066 68530
rect 186122 68474 186170 68530
rect 186226 68474 186264 68530
rect 185924 68426 186264 68474
rect 185924 68370 185962 68426
rect 186018 68370 186066 68426
rect 186122 68370 186170 68426
rect 186226 68370 186264 68426
rect 185924 68322 186264 68370
rect 185924 68266 185962 68322
rect 186018 68266 186066 68322
rect 186122 68266 186170 68322
rect 186226 68266 186264 68322
rect 185924 68238 186264 68266
rect 188768 68236 189088 69748
rect 188768 68180 188796 68236
rect 188852 68180 188900 68236
rect 188956 68180 189004 68236
rect 189060 68180 189088 68236
rect 184448 67870 184524 67898
rect 184448 67814 184458 67870
rect 184514 67814 184524 67870
rect 184448 67766 184524 67814
rect 184448 67710 184458 67766
rect 184514 67710 184524 67766
rect 184448 67662 184524 67710
rect 184448 67606 184458 67662
rect 184514 67606 184524 67662
rect 184448 67578 184524 67606
rect 185264 67870 185604 67898
rect 185264 67814 185302 67870
rect 185358 67814 185406 67870
rect 185462 67814 185510 67870
rect 185566 67814 185604 67870
rect 185264 67766 185604 67814
rect 185264 67710 185302 67766
rect 185358 67710 185406 67766
rect 185462 67710 185510 67766
rect 185566 67710 185604 67766
rect 185264 67662 185604 67710
rect 185264 67606 185302 67662
rect 185358 67606 185406 67662
rect 185462 67606 185510 67662
rect 185566 67606 185604 67662
rect 185264 67578 185604 67606
rect 188768 67870 189088 68180
rect 188768 67814 188796 67870
rect 188852 67814 188900 67870
rect 188956 67814 189004 67870
rect 189060 67814 189088 67870
rect 188768 67766 189088 67814
rect 188768 67710 188796 67766
rect 188852 67710 188900 67766
rect 188956 67710 189004 67766
rect 189060 67710 189088 67766
rect 188768 67662 189088 67710
rect 188768 67606 188796 67662
rect 188852 67606 188900 67662
rect 188956 67606 189004 67662
rect 189060 67606 189088 67662
rect 188768 66668 189088 67606
rect 188768 66612 188796 66668
rect 188852 66612 188900 66668
rect 188956 66612 189004 66668
rect 189060 66612 189088 66668
rect 188768 65100 189088 66612
rect 188768 65044 188796 65100
rect 188852 65044 188900 65100
rect 188956 65044 189004 65100
rect 189060 65044 189088 65100
rect 188768 63532 189088 65044
rect 188768 63476 188796 63532
rect 188852 63476 188900 63532
rect 188956 63476 189004 63532
rect 189060 63476 189088 63532
rect 188768 61964 189088 63476
rect 188768 61908 188796 61964
rect 188852 61908 188900 61964
rect 188956 61908 189004 61964
rect 189060 61908 189088 61964
rect 188768 60396 189088 61908
rect 188768 60340 188796 60396
rect 188852 60340 188900 60396
rect 188956 60340 189004 60396
rect 189060 60340 189088 60396
rect 188768 58828 189088 60340
rect 188768 58772 188796 58828
rect 188852 58772 188900 58828
rect 188956 58772 189004 58828
rect 189060 58772 189088 58828
rect 188768 57260 189088 58772
rect 188768 57204 188796 57260
rect 188852 57204 188900 57260
rect 188956 57204 189004 57260
rect 189060 57204 189088 57260
rect 188768 55692 189088 57204
rect 188768 55636 188796 55692
rect 188852 55636 188900 55692
rect 188956 55636 189004 55692
rect 189060 55636 189088 55692
rect 188768 54124 189088 55636
rect 188768 54068 188796 54124
rect 188852 54068 188900 54124
rect 188956 54068 189004 54124
rect 189060 54068 189088 54124
rect 188768 52556 189088 54068
rect 188768 52500 188796 52556
rect 188852 52500 188900 52556
rect 188956 52500 189004 52556
rect 189060 52500 189088 52556
rect 188768 50988 189088 52500
rect 188768 50932 188796 50988
rect 188852 50932 188900 50988
rect 188956 50932 189004 50988
rect 189060 50932 189088 50988
rect 188768 49420 189088 50932
rect 188768 49364 188796 49420
rect 188852 49364 188900 49420
rect 188956 49364 189004 49420
rect 189060 49364 189088 49420
rect 188768 47852 189088 49364
rect 188768 47796 188796 47852
rect 188852 47796 188900 47852
rect 188956 47796 189004 47852
rect 189060 47796 189088 47852
rect 188768 46284 189088 47796
rect 188768 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189088 46284
rect 188768 44716 189088 46228
rect 188768 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189088 44716
rect 188768 43148 189088 44660
rect 188768 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189088 43148
rect 188768 41580 189088 43092
rect 188768 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189088 41580
rect 188768 40012 189088 41524
rect 188768 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189088 40012
rect 188768 38444 189088 39956
rect 188768 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189088 38444
rect 158708 37838 158736 37894
rect 158792 37838 158840 37894
rect 158896 37838 158944 37894
rect 159000 37838 159028 37894
rect 158708 37790 159028 37838
rect 158708 37734 158736 37790
rect 158792 37734 158840 37790
rect 158896 37734 158944 37790
rect 159000 37734 159028 37790
rect 158708 37686 159028 37734
rect 158708 37630 158736 37686
rect 158792 37630 158840 37686
rect 158896 37630 158944 37686
rect 159000 37630 159028 37686
rect 158708 17276 159028 37630
rect 161240 37894 161316 37922
rect 161240 37838 161250 37894
rect 161306 37838 161316 37894
rect 161240 37790 161316 37838
rect 161240 37734 161250 37790
rect 161306 37734 161316 37790
rect 161240 37686 161316 37734
rect 161240 37630 161250 37686
rect 161306 37630 161316 37686
rect 161240 37602 161316 37630
rect 185924 37894 186264 37922
rect 185924 37838 185962 37894
rect 186018 37838 186066 37894
rect 186122 37838 186170 37894
rect 186226 37838 186264 37894
rect 185924 37790 186264 37838
rect 185924 37734 185962 37790
rect 186018 37734 186066 37790
rect 186122 37734 186170 37790
rect 186226 37734 186264 37790
rect 185924 37686 186264 37734
rect 185924 37630 185962 37686
rect 186018 37630 186066 37686
rect 186122 37630 186170 37686
rect 186226 37630 186264 37686
rect 185924 37602 186264 37630
rect 185264 37234 185604 37262
rect 185264 37178 185302 37234
rect 185358 37178 185406 37234
rect 185462 37178 185510 37234
rect 185566 37178 185604 37234
rect 185264 37130 185604 37178
rect 185264 37074 185302 37130
rect 185358 37074 185406 37130
rect 185462 37074 185510 37130
rect 185566 37074 185604 37130
rect 185264 37026 185604 37074
rect 185264 36970 185302 37026
rect 185358 36970 185406 37026
rect 185462 36970 185510 37026
rect 185566 36970 185604 37026
rect 185264 36942 185604 36970
rect 188768 37234 189088 38388
rect 188768 37178 188796 37234
rect 188852 37178 188900 37234
rect 188956 37178 189004 37234
rect 189060 37178 189088 37234
rect 188768 37130 189088 37178
rect 188768 37074 188796 37130
rect 188852 37074 188900 37130
rect 188956 37074 189004 37130
rect 189060 37074 189088 37130
rect 188768 37026 189088 37074
rect 188768 36970 188796 37026
rect 188852 36970 188900 37026
rect 188956 36970 189004 37026
rect 189060 36970 189088 37026
rect 158708 17220 158736 17276
rect 158792 17220 158840 17276
rect 158896 17220 158944 17276
rect 159000 17220 159028 17276
rect 158708 15708 159028 17220
rect 158708 15652 158736 15708
rect 158792 15652 158840 15708
rect 158896 15652 158944 15708
rect 159000 15652 159028 15708
rect 158708 14140 159028 15652
rect 158708 14084 158736 14140
rect 158792 14084 158840 14140
rect 158896 14084 158944 14140
rect 159000 14084 159028 14140
rect 158708 12572 159028 14084
rect 158708 12516 158736 12572
rect 158792 12516 158840 12572
rect 158896 12516 158944 12572
rect 159000 12516 159028 12572
rect 158708 11004 159028 12516
rect 158708 10948 158736 11004
rect 158792 10948 158840 11004
rect 158896 10948 158944 11004
rect 159000 10948 159028 11004
rect 158708 9436 159028 10948
rect 158708 9380 158736 9436
rect 158792 9380 158840 9436
rect 158896 9380 158944 9436
rect 159000 9380 159028 9436
rect 158708 7868 159028 9380
rect 158708 7812 158736 7868
rect 158792 7812 158840 7868
rect 158896 7812 158944 7868
rect 159000 7812 159028 7868
rect 158708 7258 159028 7812
rect 158708 7202 158736 7258
rect 158792 7202 158840 7258
rect 158896 7202 158944 7258
rect 159000 7202 159028 7258
rect 158708 7154 159028 7202
rect 158708 7098 158736 7154
rect 158792 7098 158840 7154
rect 158896 7098 158944 7154
rect 159000 7098 159028 7154
rect 158708 7050 159028 7098
rect 158708 6994 158736 7050
rect 158792 6994 158840 7050
rect 158896 6994 158944 7050
rect 159000 6994 159028 7050
rect 158708 6300 159028 6994
rect 158708 6244 158736 6300
rect 158792 6244 158840 6300
rect 158896 6244 158944 6300
rect 159000 6244 159028 6300
rect 158708 4732 159028 6244
rect 158708 4676 158736 4732
rect 158792 4676 158840 4732
rect 158896 4676 158944 4732
rect 159000 4676 159028 4732
rect 158708 3164 159028 4676
rect 158708 3108 158736 3164
rect 158792 3108 158840 3164
rect 158896 3108 158944 3164
rect 159000 3108 159028 3164
rect 158708 3076 159028 3108
rect 188768 36876 189088 36970
rect 188768 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189088 36876
rect 188768 35308 189088 36820
rect 188768 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189088 35308
rect 188768 33740 189088 35252
rect 188768 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189088 33740
rect 188768 32172 189088 33684
rect 188768 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189088 32172
rect 188768 30604 189088 32116
rect 188768 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189088 30604
rect 188768 29036 189088 30548
rect 188768 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189088 29036
rect 188768 27468 189088 28980
rect 188768 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189088 27468
rect 188768 25900 189088 27412
rect 188768 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189088 25900
rect 188768 24332 189088 25844
rect 188768 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189088 24332
rect 188768 22764 189088 24276
rect 188768 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189088 22764
rect 188768 21196 189088 22708
rect 188768 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189088 21196
rect 188768 19628 189088 21140
rect 188768 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189088 19628
rect 188768 18060 189088 19572
rect 188768 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189088 18060
rect 188768 16492 189088 18004
rect 188768 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189088 16492
rect 188768 14924 189088 16436
rect 188768 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189088 14924
rect 188768 13356 189088 14868
rect 188768 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189088 13356
rect 188768 11788 189088 13300
rect 188768 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189088 11788
rect 188768 10220 189088 11732
rect 188768 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189088 10220
rect 188768 8652 189088 10164
rect 188768 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189088 8652
rect 188768 7084 189088 8596
rect 188768 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189088 7084
rect 188768 6598 189088 7028
rect 188768 6542 188796 6598
rect 188852 6542 188900 6598
rect 188956 6542 189004 6598
rect 189060 6542 189088 6598
rect 188768 6494 189088 6542
rect 188768 6438 188796 6494
rect 188852 6438 188900 6494
rect 188956 6438 189004 6494
rect 189060 6438 189088 6494
rect 188768 6390 189088 6438
rect 188768 6334 188796 6390
rect 188852 6334 188900 6390
rect 188956 6334 189004 6390
rect 189060 6334 189088 6390
rect 188768 5516 189088 6334
rect 188768 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189088 5516
rect 188768 3948 189088 5460
rect 188768 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189088 3948
rect 188768 3076 189088 3892
rect 189428 156828 189748 156860
rect 189428 156772 189456 156828
rect 189512 156772 189560 156828
rect 189616 156772 189664 156828
rect 189720 156772 189748 156828
rect 189428 155260 189748 156772
rect 189428 155204 189456 155260
rect 189512 155204 189560 155260
rect 189616 155204 189664 155260
rect 189720 155204 189748 155260
rect 189428 153692 189748 155204
rect 189428 153636 189456 153692
rect 189512 153636 189560 153692
rect 189616 153636 189664 153692
rect 189720 153636 189748 153692
rect 189428 152124 189748 153636
rect 189428 152068 189456 152124
rect 189512 152068 189560 152124
rect 189616 152068 189664 152124
rect 189720 152068 189748 152124
rect 189428 150556 189748 152068
rect 189428 150500 189456 150556
rect 189512 150500 189560 150556
rect 189616 150500 189664 150556
rect 189720 150500 189748 150556
rect 189428 148988 189748 150500
rect 189428 148932 189456 148988
rect 189512 148932 189560 148988
rect 189616 148932 189664 148988
rect 189720 148932 189748 148988
rect 189428 147420 189748 148932
rect 189428 147364 189456 147420
rect 189512 147364 189560 147420
rect 189616 147364 189664 147420
rect 189720 147364 189748 147420
rect 189428 145852 189748 147364
rect 189428 145796 189456 145852
rect 189512 145796 189560 145852
rect 189616 145796 189664 145852
rect 189720 145796 189748 145852
rect 189428 144284 189748 145796
rect 189428 144228 189456 144284
rect 189512 144228 189560 144284
rect 189616 144228 189664 144284
rect 189720 144228 189748 144284
rect 189428 142716 189748 144228
rect 189428 142660 189456 142716
rect 189512 142660 189560 142716
rect 189616 142660 189664 142716
rect 189720 142660 189748 142716
rect 189428 141148 189748 142660
rect 189428 141092 189456 141148
rect 189512 141092 189560 141148
rect 189616 141092 189664 141148
rect 189720 141092 189748 141148
rect 189428 139580 189748 141092
rect 189428 139524 189456 139580
rect 189512 139524 189560 139580
rect 189616 139524 189664 139580
rect 189720 139524 189748 139580
rect 189428 138012 189748 139524
rect 189428 137956 189456 138012
rect 189512 137956 189560 138012
rect 189616 137956 189664 138012
rect 189720 137956 189748 138012
rect 189428 136444 189748 137956
rect 189428 136388 189456 136444
rect 189512 136388 189560 136444
rect 189616 136388 189664 136444
rect 189720 136388 189748 136444
rect 189428 134876 189748 136388
rect 189428 134820 189456 134876
rect 189512 134820 189560 134876
rect 189616 134820 189664 134876
rect 189720 134820 189748 134876
rect 189428 133308 189748 134820
rect 189428 133252 189456 133308
rect 189512 133252 189560 133308
rect 189616 133252 189664 133308
rect 189720 133252 189748 133308
rect 189428 131740 189748 133252
rect 189428 131684 189456 131740
rect 189512 131684 189560 131740
rect 189616 131684 189664 131740
rect 189720 131684 189748 131740
rect 189428 130172 189748 131684
rect 189428 130116 189456 130172
rect 189512 130116 189560 130172
rect 189616 130116 189664 130172
rect 189720 130116 189748 130172
rect 189428 129802 189748 130116
rect 189428 129746 189456 129802
rect 189512 129746 189560 129802
rect 189616 129746 189664 129802
rect 189720 129746 189748 129802
rect 189428 129698 189748 129746
rect 189428 129642 189456 129698
rect 189512 129642 189560 129698
rect 189616 129642 189664 129698
rect 189720 129642 189748 129698
rect 189428 129594 189748 129642
rect 189428 129538 189456 129594
rect 189512 129538 189560 129594
rect 189616 129538 189664 129594
rect 189720 129538 189748 129594
rect 189428 128604 189748 129538
rect 189428 128548 189456 128604
rect 189512 128548 189560 128604
rect 189616 128548 189664 128604
rect 189720 128548 189748 128604
rect 189428 127036 189748 128548
rect 189428 126980 189456 127036
rect 189512 126980 189560 127036
rect 189616 126980 189664 127036
rect 189720 126980 189748 127036
rect 189428 125468 189748 126980
rect 189428 125412 189456 125468
rect 189512 125412 189560 125468
rect 189616 125412 189664 125468
rect 189720 125412 189748 125468
rect 189428 123900 189748 125412
rect 189428 123844 189456 123900
rect 189512 123844 189560 123900
rect 189616 123844 189664 123900
rect 189720 123844 189748 123900
rect 189428 122332 189748 123844
rect 189428 122276 189456 122332
rect 189512 122276 189560 122332
rect 189616 122276 189664 122332
rect 189720 122276 189748 122332
rect 189428 120764 189748 122276
rect 189428 120708 189456 120764
rect 189512 120708 189560 120764
rect 189616 120708 189664 120764
rect 189720 120708 189748 120764
rect 189428 119196 189748 120708
rect 189428 119140 189456 119196
rect 189512 119140 189560 119196
rect 189616 119140 189664 119196
rect 189720 119140 189748 119196
rect 189428 117628 189748 119140
rect 189428 117572 189456 117628
rect 189512 117572 189560 117628
rect 189616 117572 189664 117628
rect 189720 117572 189748 117628
rect 189428 116060 189748 117572
rect 189428 116004 189456 116060
rect 189512 116004 189560 116060
rect 189616 116004 189664 116060
rect 189720 116004 189748 116060
rect 189428 114492 189748 116004
rect 189428 114436 189456 114492
rect 189512 114436 189560 114492
rect 189616 114436 189664 114492
rect 189720 114436 189748 114492
rect 189428 112924 189748 114436
rect 189428 112868 189456 112924
rect 189512 112868 189560 112924
rect 189616 112868 189664 112924
rect 189720 112868 189748 112924
rect 189428 111356 189748 112868
rect 189428 111300 189456 111356
rect 189512 111300 189560 111356
rect 189616 111300 189664 111356
rect 189720 111300 189748 111356
rect 189428 109788 189748 111300
rect 189428 109732 189456 109788
rect 189512 109732 189560 109788
rect 189616 109732 189664 109788
rect 189720 109732 189748 109788
rect 189428 108220 189748 109732
rect 189428 108164 189456 108220
rect 189512 108164 189560 108220
rect 189616 108164 189664 108220
rect 189720 108164 189748 108220
rect 189428 106652 189748 108164
rect 189428 106596 189456 106652
rect 189512 106596 189560 106652
rect 189616 106596 189664 106652
rect 189720 106596 189748 106652
rect 189428 105084 189748 106596
rect 189428 105028 189456 105084
rect 189512 105028 189560 105084
rect 189616 105028 189664 105084
rect 189720 105028 189748 105084
rect 189428 103516 189748 105028
rect 189428 103460 189456 103516
rect 189512 103460 189560 103516
rect 189616 103460 189664 103516
rect 189720 103460 189748 103516
rect 189428 101948 189748 103460
rect 189428 101892 189456 101948
rect 189512 101892 189560 101948
rect 189616 101892 189664 101948
rect 189720 101892 189748 101948
rect 189428 100380 189748 101892
rect 189428 100324 189456 100380
rect 189512 100324 189560 100380
rect 189616 100324 189664 100380
rect 189720 100324 189748 100380
rect 189428 99166 189748 100324
rect 189428 99110 189456 99166
rect 189512 99110 189560 99166
rect 189616 99110 189664 99166
rect 189720 99110 189748 99166
rect 189428 99062 189748 99110
rect 189428 99006 189456 99062
rect 189512 99006 189560 99062
rect 189616 99006 189664 99062
rect 189720 99006 189748 99062
rect 189428 98958 189748 99006
rect 189428 98902 189456 98958
rect 189512 98902 189560 98958
rect 189616 98902 189664 98958
rect 189720 98902 189748 98958
rect 189428 98812 189748 98902
rect 189428 98756 189456 98812
rect 189512 98756 189560 98812
rect 189616 98756 189664 98812
rect 189720 98756 189748 98812
rect 189428 97244 189748 98756
rect 189428 97188 189456 97244
rect 189512 97188 189560 97244
rect 189616 97188 189664 97244
rect 189720 97188 189748 97244
rect 189428 95676 189748 97188
rect 189428 95620 189456 95676
rect 189512 95620 189560 95676
rect 189616 95620 189664 95676
rect 189720 95620 189748 95676
rect 189428 94108 189748 95620
rect 189428 94052 189456 94108
rect 189512 94052 189560 94108
rect 189616 94052 189664 94108
rect 189720 94052 189748 94108
rect 189428 92540 189748 94052
rect 189428 92484 189456 92540
rect 189512 92484 189560 92540
rect 189616 92484 189664 92540
rect 189720 92484 189748 92540
rect 189428 90972 189748 92484
rect 189428 90916 189456 90972
rect 189512 90916 189560 90972
rect 189616 90916 189664 90972
rect 189720 90916 189748 90972
rect 189428 89404 189748 90916
rect 189428 89348 189456 89404
rect 189512 89348 189560 89404
rect 189616 89348 189664 89404
rect 189720 89348 189748 89404
rect 189428 87836 189748 89348
rect 189428 87780 189456 87836
rect 189512 87780 189560 87836
rect 189616 87780 189664 87836
rect 189720 87780 189748 87836
rect 189428 86268 189748 87780
rect 189428 86212 189456 86268
rect 189512 86212 189560 86268
rect 189616 86212 189664 86268
rect 189720 86212 189748 86268
rect 189428 84700 189748 86212
rect 189428 84644 189456 84700
rect 189512 84644 189560 84700
rect 189616 84644 189664 84700
rect 189720 84644 189748 84700
rect 189428 83132 189748 84644
rect 189428 83076 189456 83132
rect 189512 83076 189560 83132
rect 189616 83076 189664 83132
rect 189720 83076 189748 83132
rect 189428 81564 189748 83076
rect 189428 81508 189456 81564
rect 189512 81508 189560 81564
rect 189616 81508 189664 81564
rect 189720 81508 189748 81564
rect 189428 79996 189748 81508
rect 189428 79940 189456 79996
rect 189512 79940 189560 79996
rect 189616 79940 189664 79996
rect 189720 79940 189748 79996
rect 189428 78428 189748 79940
rect 189428 78372 189456 78428
rect 189512 78372 189560 78428
rect 189616 78372 189664 78428
rect 189720 78372 189748 78428
rect 189428 76860 189748 78372
rect 189428 76804 189456 76860
rect 189512 76804 189560 76860
rect 189616 76804 189664 76860
rect 189720 76804 189748 76860
rect 189428 75292 189748 76804
rect 189428 75236 189456 75292
rect 189512 75236 189560 75292
rect 189616 75236 189664 75292
rect 189720 75236 189748 75292
rect 189428 73724 189748 75236
rect 189428 73668 189456 73724
rect 189512 73668 189560 73724
rect 189616 73668 189664 73724
rect 189720 73668 189748 73724
rect 189428 72156 189748 73668
rect 189428 72100 189456 72156
rect 189512 72100 189560 72156
rect 189616 72100 189664 72156
rect 189720 72100 189748 72156
rect 189428 70588 189748 72100
rect 189428 70532 189456 70588
rect 189512 70532 189560 70588
rect 189616 70532 189664 70588
rect 189720 70532 189748 70588
rect 189428 69020 189748 70532
rect 189428 68964 189456 69020
rect 189512 68964 189560 69020
rect 189616 68964 189664 69020
rect 189720 68964 189748 69020
rect 189428 68530 189748 68964
rect 189428 68474 189456 68530
rect 189512 68474 189560 68530
rect 189616 68474 189664 68530
rect 189720 68474 189748 68530
rect 189428 68426 189748 68474
rect 189428 68370 189456 68426
rect 189512 68370 189560 68426
rect 189616 68370 189664 68426
rect 189720 68370 189748 68426
rect 189428 68322 189748 68370
rect 189428 68266 189456 68322
rect 189512 68266 189560 68322
rect 189616 68266 189664 68322
rect 189720 68266 189748 68322
rect 189428 67452 189748 68266
rect 189428 67396 189456 67452
rect 189512 67396 189560 67452
rect 189616 67396 189664 67452
rect 189720 67396 189748 67452
rect 189428 65884 189748 67396
rect 189428 65828 189456 65884
rect 189512 65828 189560 65884
rect 189616 65828 189664 65884
rect 189720 65828 189748 65884
rect 189428 64316 189748 65828
rect 189428 64260 189456 64316
rect 189512 64260 189560 64316
rect 189616 64260 189664 64316
rect 189720 64260 189748 64316
rect 189428 62748 189748 64260
rect 189428 62692 189456 62748
rect 189512 62692 189560 62748
rect 189616 62692 189664 62748
rect 189720 62692 189748 62748
rect 189428 61180 189748 62692
rect 189428 61124 189456 61180
rect 189512 61124 189560 61180
rect 189616 61124 189664 61180
rect 189720 61124 189748 61180
rect 189428 59612 189748 61124
rect 189428 59556 189456 59612
rect 189512 59556 189560 59612
rect 189616 59556 189664 59612
rect 189720 59556 189748 59612
rect 189428 58044 189748 59556
rect 189428 57988 189456 58044
rect 189512 57988 189560 58044
rect 189616 57988 189664 58044
rect 189720 57988 189748 58044
rect 189428 56476 189748 57988
rect 189428 56420 189456 56476
rect 189512 56420 189560 56476
rect 189616 56420 189664 56476
rect 189720 56420 189748 56476
rect 189428 54908 189748 56420
rect 189428 54852 189456 54908
rect 189512 54852 189560 54908
rect 189616 54852 189664 54908
rect 189720 54852 189748 54908
rect 189428 53340 189748 54852
rect 189428 53284 189456 53340
rect 189512 53284 189560 53340
rect 189616 53284 189664 53340
rect 189720 53284 189748 53340
rect 189428 51772 189748 53284
rect 189428 51716 189456 51772
rect 189512 51716 189560 51772
rect 189616 51716 189664 51772
rect 189720 51716 189748 51772
rect 189428 50204 189748 51716
rect 189428 50148 189456 50204
rect 189512 50148 189560 50204
rect 189616 50148 189664 50204
rect 189720 50148 189748 50204
rect 189428 48636 189748 50148
rect 189428 48580 189456 48636
rect 189512 48580 189560 48636
rect 189616 48580 189664 48636
rect 189720 48580 189748 48636
rect 189428 47068 189748 48580
rect 189428 47012 189456 47068
rect 189512 47012 189560 47068
rect 189616 47012 189664 47068
rect 189720 47012 189748 47068
rect 189428 45500 189748 47012
rect 189428 45444 189456 45500
rect 189512 45444 189560 45500
rect 189616 45444 189664 45500
rect 189720 45444 189748 45500
rect 189428 43932 189748 45444
rect 189428 43876 189456 43932
rect 189512 43876 189560 43932
rect 189616 43876 189664 43932
rect 189720 43876 189748 43932
rect 189428 42364 189748 43876
rect 189428 42308 189456 42364
rect 189512 42308 189560 42364
rect 189616 42308 189664 42364
rect 189720 42308 189748 42364
rect 189428 40796 189748 42308
rect 189428 40740 189456 40796
rect 189512 40740 189560 40796
rect 189616 40740 189664 40796
rect 189720 40740 189748 40796
rect 189428 39228 189748 40740
rect 189428 39172 189456 39228
rect 189512 39172 189560 39228
rect 189616 39172 189664 39228
rect 189720 39172 189748 39228
rect 189428 37894 189748 39172
rect 189428 37838 189456 37894
rect 189512 37838 189560 37894
rect 189616 37838 189664 37894
rect 189720 37838 189748 37894
rect 189428 37790 189748 37838
rect 189428 37734 189456 37790
rect 189512 37734 189560 37790
rect 189616 37734 189664 37790
rect 189720 37734 189748 37790
rect 189428 37686 189748 37734
rect 189428 37604 189456 37686
rect 189512 37604 189560 37686
rect 189616 37604 189664 37686
rect 189720 37604 189748 37686
rect 189428 36092 189748 37604
rect 189428 36036 189456 36092
rect 189512 36036 189560 36092
rect 189616 36036 189664 36092
rect 189720 36036 189748 36092
rect 189428 34524 189748 36036
rect 189428 34468 189456 34524
rect 189512 34468 189560 34524
rect 189616 34468 189664 34524
rect 189720 34468 189748 34524
rect 189428 32956 189748 34468
rect 189428 32900 189456 32956
rect 189512 32900 189560 32956
rect 189616 32900 189664 32956
rect 189720 32900 189748 32956
rect 189428 31388 189748 32900
rect 189428 31332 189456 31388
rect 189512 31332 189560 31388
rect 189616 31332 189664 31388
rect 189720 31332 189748 31388
rect 189428 29820 189748 31332
rect 189428 29764 189456 29820
rect 189512 29764 189560 29820
rect 189616 29764 189664 29820
rect 189720 29764 189748 29820
rect 189428 28252 189748 29764
rect 189428 28196 189456 28252
rect 189512 28196 189560 28252
rect 189616 28196 189664 28252
rect 189720 28196 189748 28252
rect 189428 26684 189748 28196
rect 189428 26628 189456 26684
rect 189512 26628 189560 26684
rect 189616 26628 189664 26684
rect 189720 26628 189748 26684
rect 189428 25116 189748 26628
rect 189428 25060 189456 25116
rect 189512 25060 189560 25116
rect 189616 25060 189664 25116
rect 189720 25060 189748 25116
rect 189428 23548 189748 25060
rect 189428 23492 189456 23548
rect 189512 23492 189560 23548
rect 189616 23492 189664 23548
rect 189720 23492 189748 23548
rect 189428 21980 189748 23492
rect 189428 21924 189456 21980
rect 189512 21924 189560 21980
rect 189616 21924 189664 21980
rect 189720 21924 189748 21980
rect 189428 20412 189748 21924
rect 189428 20356 189456 20412
rect 189512 20356 189560 20412
rect 189616 20356 189664 20412
rect 189720 20356 189748 20412
rect 189428 18844 189748 20356
rect 189428 18788 189456 18844
rect 189512 18788 189560 18844
rect 189616 18788 189664 18844
rect 189720 18788 189748 18844
rect 189428 17276 189748 18788
rect 189428 17220 189456 17276
rect 189512 17220 189560 17276
rect 189616 17220 189664 17276
rect 189720 17220 189748 17276
rect 189428 15708 189748 17220
rect 189428 15652 189456 15708
rect 189512 15652 189560 15708
rect 189616 15652 189664 15708
rect 189720 15652 189748 15708
rect 189428 14140 189748 15652
rect 189428 14084 189456 14140
rect 189512 14084 189560 14140
rect 189616 14084 189664 14140
rect 189720 14084 189748 14140
rect 189428 12572 189748 14084
rect 189428 12516 189456 12572
rect 189512 12516 189560 12572
rect 189616 12516 189664 12572
rect 189720 12516 189748 12572
rect 189428 11004 189748 12516
rect 189428 10948 189456 11004
rect 189512 10948 189560 11004
rect 189616 10948 189664 11004
rect 189720 10948 189748 11004
rect 189428 9436 189748 10948
rect 189428 9380 189456 9436
rect 189512 9380 189560 9436
rect 189616 9380 189664 9436
rect 189720 9380 189748 9436
rect 189428 7868 189748 9380
rect 189428 7812 189456 7868
rect 189512 7812 189560 7868
rect 189616 7812 189664 7868
rect 189720 7812 189748 7868
rect 189428 7258 189748 7812
rect 189428 7202 189456 7258
rect 189512 7202 189560 7258
rect 189616 7202 189664 7258
rect 189720 7202 189748 7258
rect 189428 7154 189748 7202
rect 189428 7098 189456 7154
rect 189512 7098 189560 7154
rect 189616 7098 189664 7154
rect 189720 7098 189748 7154
rect 189428 7050 189748 7098
rect 189428 6994 189456 7050
rect 189512 6994 189560 7050
rect 189616 6994 189664 7050
rect 189720 6994 189748 7050
rect 189428 6300 189748 6994
rect 189428 6244 189456 6300
rect 189512 6244 189560 6300
rect 189616 6244 189664 6300
rect 189720 6244 189748 6300
rect 189428 4732 189748 6244
rect 189428 4676 189456 4732
rect 189512 4676 189560 4732
rect 189616 4676 189664 4732
rect 189720 4676 189748 4732
rect 189428 3164 189748 4676
rect 189428 3108 189456 3164
rect 189512 3108 189560 3164
rect 189616 3108 189664 3164
rect 189720 3108 189748 3164
rect 189428 3076 189748 3108
<< via4 >>
rect 4476 129086 4532 129142
rect 4580 129086 4636 129142
rect 4684 129086 4740 129142
rect 4476 128982 4532 129038
rect 4580 128982 4636 129038
rect 4684 128982 4740 129038
rect 4476 128878 4532 128934
rect 4580 128878 4636 128934
rect 4684 128878 4740 128934
rect 4476 98450 4532 98506
rect 4580 98450 4636 98506
rect 4684 98450 4740 98506
rect 4476 98346 4532 98402
rect 4580 98346 4636 98402
rect 4684 98346 4740 98402
rect 4476 98242 4532 98298
rect 4580 98242 4636 98298
rect 4684 98242 4740 98298
rect 4476 67814 4532 67870
rect 4580 67814 4636 67870
rect 4684 67814 4740 67870
rect 4476 67710 4532 67766
rect 4580 67710 4636 67766
rect 4684 67710 4740 67766
rect 4476 67606 4532 67662
rect 4580 67606 4636 67662
rect 4684 67606 4740 67662
rect 4476 37178 4532 37234
rect 4580 37178 4636 37234
rect 4684 37178 4740 37234
rect 4476 37074 4532 37130
rect 4580 37074 4636 37130
rect 4684 37074 4740 37130
rect 4476 36970 4532 37026
rect 4580 36970 4636 37026
rect 4684 36970 4740 37026
rect 4476 6542 4532 6598
rect 4580 6542 4636 6598
rect 4684 6542 4740 6598
rect 4476 6438 4532 6494
rect 4580 6438 4636 6494
rect 4684 6438 4740 6494
rect 4476 6334 4532 6390
rect 4580 6334 4636 6390
rect 4684 6334 4740 6390
rect 5136 129746 5192 129802
rect 5240 129746 5296 129802
rect 5344 129746 5400 129802
rect 5136 129642 5192 129698
rect 5240 129642 5296 129698
rect 5344 129642 5400 129698
rect 5136 129538 5192 129594
rect 5240 129538 5296 129594
rect 5344 129538 5400 129594
rect 20038 129746 20094 129802
rect 20142 129746 20198 129802
rect 20246 129746 20302 129802
rect 20038 129642 20094 129698
rect 20142 129642 20198 129698
rect 20246 129642 20302 129698
rect 20038 129538 20094 129594
rect 20142 129538 20198 129594
rect 20246 129538 20302 129594
rect 20698 129086 20754 129142
rect 20802 129086 20858 129142
rect 20906 129086 20962 129142
rect 20698 128982 20754 129038
rect 20802 128982 20858 129038
rect 20906 128982 20962 129038
rect 20698 128878 20754 128934
rect 20802 128878 20858 128934
rect 20906 128878 20962 128934
rect 35196 129086 35252 129142
rect 35300 129086 35356 129142
rect 35404 129086 35460 129142
rect 35196 128982 35252 129038
rect 35300 128982 35356 129038
rect 35404 128982 35460 129038
rect 35196 128878 35252 128934
rect 35300 128878 35356 128934
rect 35404 128878 35460 128934
rect 5136 99110 5192 99166
rect 5240 99110 5296 99166
rect 5344 99110 5400 99166
rect 5136 99006 5192 99062
rect 5240 99006 5296 99062
rect 5344 99006 5400 99062
rect 5136 98902 5192 98958
rect 5240 98902 5296 98958
rect 5344 98902 5400 98958
rect 20038 99110 20094 99166
rect 20142 99110 20198 99166
rect 20246 99110 20302 99166
rect 20038 99006 20094 99062
rect 20142 99006 20198 99062
rect 20246 99006 20302 99062
rect 20038 98902 20094 98958
rect 20142 98902 20198 98958
rect 20246 98902 20302 98958
rect 20698 98450 20754 98506
rect 20802 98450 20858 98506
rect 20906 98450 20962 98506
rect 20698 98346 20754 98402
rect 20802 98346 20858 98402
rect 20906 98346 20962 98402
rect 20698 98242 20754 98298
rect 20802 98242 20858 98298
rect 20906 98242 20962 98298
rect 35196 98450 35252 98506
rect 35300 98450 35356 98506
rect 35404 98450 35460 98506
rect 35196 98346 35252 98402
rect 35300 98346 35356 98402
rect 35404 98346 35460 98402
rect 35196 98242 35252 98298
rect 35300 98242 35356 98298
rect 35404 98242 35460 98298
rect 5136 68474 5192 68530
rect 5240 68474 5296 68530
rect 5344 68474 5400 68530
rect 5136 68370 5192 68426
rect 5240 68370 5296 68426
rect 5344 68370 5400 68426
rect 5136 68266 5192 68322
rect 5240 68266 5296 68322
rect 5344 68266 5400 68322
rect 20038 68474 20094 68530
rect 20142 68474 20198 68530
rect 20246 68474 20302 68530
rect 20038 68370 20094 68426
rect 20142 68370 20198 68426
rect 20246 68370 20302 68426
rect 20038 68266 20094 68322
rect 20142 68266 20198 68322
rect 20246 68266 20302 68322
rect 20698 67814 20754 67870
rect 20802 67814 20858 67870
rect 20906 67814 20962 67870
rect 20698 67710 20754 67766
rect 20802 67710 20858 67766
rect 20906 67710 20962 67766
rect 20698 67606 20754 67662
rect 20802 67606 20858 67662
rect 20906 67606 20962 67662
rect 35196 67814 35252 67870
rect 35300 67814 35356 67870
rect 35404 67814 35460 67870
rect 35196 67710 35252 67766
rect 35300 67710 35356 67766
rect 35404 67710 35460 67766
rect 35196 67606 35252 67662
rect 35300 67606 35356 67662
rect 35404 67606 35460 67662
rect 5136 37838 5192 37894
rect 5240 37838 5296 37894
rect 5344 37838 5400 37894
rect 5136 37734 5192 37790
rect 5240 37734 5296 37790
rect 5344 37734 5400 37790
rect 5136 37660 5192 37686
rect 5136 37630 5192 37660
rect 5240 37660 5296 37686
rect 5240 37630 5296 37660
rect 5344 37660 5400 37686
rect 5344 37630 5400 37660
rect 20038 37838 20094 37894
rect 20142 37838 20198 37894
rect 20246 37838 20302 37894
rect 20038 37734 20094 37790
rect 20142 37734 20198 37790
rect 20246 37734 20302 37790
rect 20038 37630 20094 37686
rect 20142 37630 20198 37686
rect 20246 37630 20302 37686
rect 29062 37838 29118 37894
rect 29062 37734 29118 37790
rect 29062 37630 29118 37686
rect 20698 37178 20754 37234
rect 20802 37178 20858 37234
rect 20906 37178 20962 37234
rect 20698 37074 20754 37130
rect 20802 37074 20858 37130
rect 20906 37074 20962 37130
rect 20698 36970 20754 37026
rect 20802 36970 20858 37026
rect 20906 36970 20962 37026
rect 35196 37178 35252 37234
rect 35300 37178 35356 37234
rect 35404 37178 35460 37234
rect 35196 37074 35252 37130
rect 35300 37074 35356 37130
rect 35404 37074 35460 37130
rect 35196 36970 35252 37026
rect 35300 36970 35356 37026
rect 35404 36970 35460 37026
rect 5136 7202 5192 7258
rect 5240 7202 5296 7258
rect 5344 7202 5400 7258
rect 5136 7098 5192 7154
rect 5240 7098 5296 7154
rect 5344 7098 5400 7154
rect 5136 6994 5192 7050
rect 5240 6994 5296 7050
rect 5344 6994 5400 7050
rect 35196 6542 35252 6598
rect 35300 6542 35356 6598
rect 35404 6542 35460 6598
rect 35196 6438 35252 6494
rect 35300 6438 35356 6494
rect 35404 6438 35460 6494
rect 35196 6334 35252 6390
rect 35300 6334 35356 6390
rect 35404 6334 35460 6390
rect 35856 129746 35912 129802
rect 35960 129746 36016 129802
rect 36064 129746 36120 129802
rect 35856 129642 35912 129698
rect 35960 129642 36016 129698
rect 36064 129642 36120 129698
rect 35856 129538 35912 129594
rect 35960 129538 36016 129594
rect 36064 129538 36120 129594
rect 48528 129746 48584 129802
rect 48528 129642 48584 129698
rect 48528 129538 48584 129594
rect 49962 129746 50018 129802
rect 49962 129642 50018 129698
rect 49962 129538 50018 129594
rect 51414 129746 51470 129802
rect 51414 129642 51470 129698
rect 51414 129538 51470 129594
rect 54666 129746 54722 129802
rect 54666 129642 54722 129698
rect 54666 129538 54722 129594
rect 65732 129746 65788 129802
rect 65732 129642 65788 129698
rect 65732 129538 65788 129594
rect 66576 129746 66632 129802
rect 66680 129746 66736 129802
rect 66784 129746 66840 129802
rect 66576 129642 66632 129698
rect 66680 129642 66736 129698
rect 66784 129642 66840 129698
rect 66576 129538 66632 129594
rect 66680 129538 66736 129594
rect 66784 129538 66840 129594
rect 49598 129086 49654 129142
rect 49598 128982 49654 129038
rect 49598 128878 49654 128934
rect 50598 129086 50654 129142
rect 50598 128982 50654 129038
rect 50598 128878 50654 128934
rect 52039 129086 52095 129142
rect 52039 128982 52095 129038
rect 52039 128878 52095 128934
rect 60826 129086 60882 129142
rect 60826 128982 60882 129038
rect 60826 128878 60882 128934
rect 65296 129086 65352 129142
rect 65296 128982 65352 129038
rect 65296 128878 65352 128934
rect 35856 99110 35912 99166
rect 35960 99110 36016 99166
rect 36064 99110 36120 99166
rect 35856 99006 35912 99062
rect 35960 99006 36016 99062
rect 36064 99006 36120 99062
rect 35856 98902 35912 98958
rect 35960 98902 36016 98958
rect 36064 98902 36120 98958
rect 48528 99110 48584 99166
rect 48528 99006 48584 99062
rect 48528 98902 48584 98958
rect 49962 99110 50018 99166
rect 49962 99006 50018 99062
rect 49962 98902 50018 98958
rect 51414 99110 51470 99166
rect 51414 99006 51470 99062
rect 51414 98902 51470 98958
rect 54666 99110 54722 99166
rect 54666 99006 54722 99062
rect 54666 98902 54722 98958
rect 65732 99110 65788 99166
rect 65732 99006 65788 99062
rect 65732 98902 65788 98958
rect 66576 99110 66632 99166
rect 66680 99110 66736 99166
rect 66784 99110 66840 99166
rect 66576 99006 66632 99062
rect 66680 99006 66736 99062
rect 66784 99006 66840 99062
rect 66576 98902 66632 98958
rect 66680 98902 66736 98958
rect 66784 98902 66840 98958
rect 49598 98450 49654 98506
rect 49598 98346 49654 98402
rect 49598 98242 49654 98298
rect 50598 98450 50654 98506
rect 50598 98346 50654 98402
rect 50598 98242 50654 98298
rect 52039 98450 52095 98506
rect 52039 98346 52095 98402
rect 52039 98242 52095 98298
rect 60826 98450 60882 98506
rect 60826 98346 60882 98402
rect 60826 98242 60882 98298
rect 65296 98450 65352 98506
rect 65296 98346 65352 98402
rect 65296 98242 65352 98298
rect 35856 68474 35912 68530
rect 35960 68474 36016 68530
rect 36064 68474 36120 68530
rect 35856 68370 35912 68426
rect 35960 68370 36016 68426
rect 36064 68370 36120 68426
rect 44562 68403 44618 68459
rect 35856 68266 35912 68322
rect 35960 68266 36016 68322
rect 36064 68266 36120 68322
rect 42582 68285 42638 68341
rect 44562 68299 44618 68355
rect 48528 68474 48584 68530
rect 48528 68370 48584 68426
rect 48528 68266 48584 68322
rect 49962 68474 50018 68530
rect 49962 68370 50018 68426
rect 49962 68266 50018 68322
rect 51414 68474 51470 68530
rect 51414 68370 51470 68426
rect 51414 68266 51470 68322
rect 54666 68474 54722 68530
rect 54666 68370 54722 68426
rect 54666 68266 54722 68322
rect 65732 68474 65788 68530
rect 65732 68370 65788 68426
rect 65732 68266 65788 68322
rect 66576 68474 66632 68530
rect 66680 68474 66736 68530
rect 66784 68474 66840 68530
rect 66576 68370 66632 68426
rect 66680 68370 66736 68426
rect 66784 68370 66840 68426
rect 66576 68266 66632 68322
rect 66680 68266 66736 68322
rect 66784 68266 66840 68322
rect 44694 67799 44750 67855
rect 44694 67695 44750 67751
rect 46014 67799 46070 67855
rect 46014 67695 46070 67751
rect 49598 67814 49654 67870
rect 49598 67710 49654 67766
rect 49598 67606 49654 67662
rect 50598 67814 50654 67870
rect 50598 67710 50654 67766
rect 50598 67606 50654 67662
rect 52039 67814 52095 67870
rect 52039 67710 52095 67766
rect 52039 67606 52095 67662
rect 60826 67814 60882 67870
rect 60826 67710 60882 67766
rect 60826 67606 60882 67662
rect 65296 67814 65352 67870
rect 65296 67710 65352 67766
rect 65296 67606 65352 67662
rect 35856 37838 35912 37894
rect 35960 37838 36016 37894
rect 36064 37838 36120 37894
rect 35856 37734 35912 37790
rect 35960 37734 36016 37790
rect 36064 37734 36120 37790
rect 35856 37630 35912 37686
rect 35960 37630 36016 37686
rect 36064 37630 36120 37686
rect 43728 37838 43784 37894
rect 43728 37734 43784 37790
rect 43728 37630 43784 37686
rect 45970 37838 46026 37894
rect 45970 37734 46026 37790
rect 45970 37630 46026 37686
rect 47652 37838 47708 37894
rect 47652 37734 47708 37790
rect 47652 37630 47708 37686
rect 96636 129086 96692 129142
rect 96740 129086 96796 129142
rect 96844 129086 96900 129142
rect 96636 128982 96692 129038
rect 96740 128982 96796 129038
rect 96844 128982 96900 129038
rect 96636 128878 96692 128934
rect 96740 128878 96796 128934
rect 96844 128878 96900 128934
rect 96636 98450 96692 98506
rect 96740 98450 96796 98506
rect 96844 98450 96900 98506
rect 96636 98346 96692 98402
rect 96740 98346 96796 98402
rect 96844 98346 96900 98402
rect 96636 98242 96692 98298
rect 96740 98242 96796 98298
rect 96844 98242 96900 98298
rect 96636 67814 96692 67870
rect 96740 67814 96796 67870
rect 96844 67814 96900 67870
rect 96636 67710 96692 67766
rect 96740 67710 96796 67766
rect 96844 67710 96900 67766
rect 96636 67606 96692 67662
rect 96740 67606 96796 67662
rect 96844 67606 96900 67662
rect 97296 129746 97352 129802
rect 97400 129746 97456 129802
rect 97504 129746 97560 129802
rect 97296 129642 97352 129698
rect 97400 129642 97456 129698
rect 97504 129642 97560 129698
rect 97296 129538 97352 129594
rect 97400 129538 97456 129594
rect 97504 129538 97560 129594
rect 97296 99110 97352 99166
rect 97400 99110 97456 99166
rect 97504 99110 97560 99166
rect 97296 99006 97352 99062
rect 97400 99006 97456 99062
rect 97504 99006 97560 99062
rect 97296 98902 97352 98958
rect 97400 98902 97456 98958
rect 97504 98902 97560 98958
rect 97296 68474 97352 68530
rect 97400 68474 97456 68530
rect 97504 68474 97560 68530
rect 97296 68370 97352 68426
rect 97400 68370 97456 68426
rect 97504 68370 97560 68426
rect 97296 68266 97352 68322
rect 97400 68266 97456 68322
rect 97504 68266 97560 68322
rect 66576 37838 66632 37894
rect 66680 37838 66736 37894
rect 66784 37838 66840 37894
rect 66576 37734 66632 37790
rect 66680 37734 66736 37790
rect 66784 37734 66840 37790
rect 66576 37630 66632 37686
rect 66680 37630 66736 37686
rect 66784 37630 66840 37686
rect 40074 37178 40130 37234
rect 40074 37074 40130 37130
rect 40074 36970 40130 37026
rect 44384 37178 44440 37234
rect 44384 37074 44440 37130
rect 44384 36970 44440 37026
rect 47294 37178 47350 37234
rect 47294 37074 47350 37130
rect 47294 36970 47350 37026
rect 48308 37178 48364 37234
rect 48308 37074 48364 37130
rect 48308 36970 48364 37026
rect 97296 37838 97352 37894
rect 97400 37838 97456 37894
rect 97504 37838 97560 37894
rect 97296 37734 97352 37790
rect 97400 37734 97456 37790
rect 97504 37734 97560 37790
rect 97296 37630 97352 37686
rect 97400 37630 97456 37686
rect 97504 37630 97560 37686
rect 127356 129086 127412 129142
rect 127460 129086 127516 129142
rect 127564 129086 127620 129142
rect 127356 128982 127412 129038
rect 127460 128982 127516 129038
rect 127564 128982 127620 129038
rect 127356 128878 127412 128934
rect 127460 128878 127516 128934
rect 127564 128878 127620 128934
rect 127356 98450 127412 98506
rect 127460 98450 127516 98506
rect 127564 98450 127620 98506
rect 127356 98346 127412 98402
rect 127460 98346 127516 98402
rect 127564 98346 127620 98402
rect 127356 98242 127412 98298
rect 127460 98242 127516 98298
rect 127564 98242 127620 98298
rect 127356 67814 127412 67870
rect 127460 67814 127516 67870
rect 127564 67814 127620 67870
rect 127356 67710 127412 67766
rect 127460 67710 127516 67766
rect 127564 67710 127620 67766
rect 127356 67606 127412 67662
rect 127460 67606 127516 67662
rect 127564 67606 127620 67662
rect 127356 37178 127412 37234
rect 127460 37178 127516 37234
rect 127564 37178 127620 37234
rect 127356 37074 127412 37130
rect 127460 37074 127516 37130
rect 127564 37074 127620 37130
rect 127356 36970 127412 37026
rect 127460 36970 127516 37026
rect 127564 36970 127620 37026
rect 128016 129746 128072 129802
rect 128120 129746 128176 129802
rect 128224 129746 128280 129802
rect 128016 129642 128072 129698
rect 128120 129642 128176 129698
rect 128224 129642 128280 129698
rect 128016 129538 128072 129594
rect 128120 129538 128176 129594
rect 128224 129538 128280 129594
rect 128016 99110 128072 99166
rect 128120 99110 128176 99166
rect 128224 99110 128280 99166
rect 128016 99006 128072 99062
rect 128120 99006 128176 99062
rect 128224 99006 128280 99062
rect 128016 98902 128072 98958
rect 128120 98902 128176 98958
rect 128224 98902 128280 98958
rect 128016 68474 128072 68530
rect 128120 68474 128176 68530
rect 128224 68474 128280 68530
rect 128016 68370 128072 68426
rect 128120 68370 128176 68426
rect 128224 68370 128280 68426
rect 128016 68266 128072 68322
rect 128120 68266 128176 68322
rect 128224 68266 128280 68322
rect 158076 129086 158132 129142
rect 158180 129086 158236 129142
rect 158284 129086 158340 129142
rect 158076 128982 158132 129038
rect 158180 128982 158236 129038
rect 158284 128982 158340 129038
rect 158076 128878 158132 128934
rect 158180 128878 158236 128934
rect 158284 128878 158340 128934
rect 158076 98450 158132 98506
rect 158180 98450 158236 98506
rect 158284 98450 158340 98506
rect 158076 98346 158132 98402
rect 158180 98346 158236 98402
rect 158284 98346 158340 98402
rect 158076 98242 158132 98298
rect 158180 98242 158236 98298
rect 158284 98242 158340 98298
rect 158076 67814 158132 67870
rect 158180 67814 158236 67870
rect 158284 67814 158340 67870
rect 158076 67710 158132 67766
rect 158180 67710 158236 67766
rect 158284 67710 158340 67766
rect 158076 67606 158132 67662
rect 158180 67606 158236 67662
rect 158284 67606 158340 67662
rect 128016 37838 128072 37894
rect 128120 37838 128176 37894
rect 128224 37838 128280 37894
rect 128016 37734 128072 37790
rect 128120 37734 128176 37790
rect 128224 37734 128280 37790
rect 128016 37630 128072 37686
rect 128120 37630 128176 37686
rect 128224 37630 128280 37686
rect 35856 7202 35912 7258
rect 35960 7202 36016 7258
rect 36064 7202 36120 7258
rect 35856 7098 35912 7154
rect 35960 7098 36016 7154
rect 36064 7098 36120 7154
rect 35856 6994 35912 7050
rect 35960 6994 36016 7050
rect 36064 6994 36120 7050
rect 65916 6542 65972 6598
rect 66020 6542 66076 6598
rect 66124 6542 66180 6598
rect 65916 6438 65972 6494
rect 66020 6438 66076 6494
rect 66124 6438 66180 6494
rect 65916 6334 65972 6390
rect 66020 6334 66076 6390
rect 66124 6334 66180 6390
rect 66576 7202 66632 7258
rect 66680 7202 66736 7258
rect 66784 7202 66840 7258
rect 66576 7098 66632 7154
rect 66680 7098 66736 7154
rect 66784 7098 66840 7154
rect 66576 6994 66632 7050
rect 66680 6994 66736 7050
rect 66784 6994 66840 7050
rect 96636 6542 96692 6598
rect 96740 6542 96796 6598
rect 96844 6542 96900 6598
rect 96636 6438 96692 6494
rect 96740 6438 96796 6494
rect 96844 6438 96900 6494
rect 96636 6334 96692 6390
rect 96740 6334 96796 6390
rect 96844 6334 96900 6390
rect 97296 7202 97352 7258
rect 97400 7202 97456 7258
rect 97504 7202 97560 7258
rect 97296 7098 97352 7154
rect 97400 7098 97456 7154
rect 97504 7098 97560 7154
rect 97296 6994 97352 7050
rect 97400 6994 97456 7050
rect 97504 6994 97560 7050
rect 127356 6542 127412 6598
rect 127460 6542 127516 6598
rect 127564 6542 127620 6598
rect 127356 6438 127412 6494
rect 127460 6438 127516 6494
rect 127564 6438 127620 6494
rect 127356 6334 127412 6390
rect 127460 6334 127516 6390
rect 127564 6334 127620 6390
rect 130890 37178 130946 37234
rect 130890 37074 130946 37130
rect 130890 36970 130946 37026
rect 158076 37178 158132 37234
rect 158180 37178 158236 37234
rect 158284 37178 158340 37234
rect 158076 37074 158132 37130
rect 158180 37074 158236 37130
rect 158284 37074 158340 37130
rect 158076 36970 158132 37026
rect 158180 36970 158236 37026
rect 158284 36970 158340 37026
rect 128016 7202 128072 7258
rect 128120 7202 128176 7258
rect 128224 7202 128280 7258
rect 128016 7098 128072 7154
rect 128120 7098 128176 7154
rect 128224 7098 128280 7154
rect 128016 6994 128072 7050
rect 128120 6994 128176 7050
rect 128224 6994 128280 7050
rect 158076 6542 158132 6598
rect 158180 6542 158236 6598
rect 158284 6542 158340 6598
rect 158076 6438 158132 6494
rect 158180 6438 158236 6494
rect 158284 6438 158340 6494
rect 158076 6334 158132 6390
rect 158180 6334 158236 6390
rect 158284 6334 158340 6390
rect 158736 129746 158792 129802
rect 158840 129746 158896 129802
rect 158944 129746 159000 129802
rect 158736 129642 158792 129698
rect 158840 129642 158896 129698
rect 158944 129642 159000 129698
rect 158736 129538 158792 129594
rect 158840 129538 158896 129594
rect 158944 129538 159000 129594
rect 184022 129746 184078 129802
rect 184022 129642 184078 129698
rect 184022 129538 184078 129594
rect 185962 129746 186018 129802
rect 186066 129746 186122 129802
rect 186170 129746 186226 129802
rect 185962 129642 186018 129698
rect 186066 129642 186122 129698
rect 186170 129642 186226 129698
rect 185962 129538 186018 129594
rect 186066 129538 186122 129594
rect 186170 129538 186226 129594
rect 184458 129086 184514 129142
rect 184458 128982 184514 129038
rect 184458 128878 184514 128934
rect 185302 129086 185358 129142
rect 185406 129086 185462 129142
rect 185510 129086 185566 129142
rect 185302 128982 185358 129038
rect 185406 128982 185462 129038
rect 185510 128982 185566 129038
rect 185302 128878 185358 128934
rect 185406 128878 185462 128934
rect 185510 128878 185566 128934
rect 188796 129086 188852 129142
rect 188900 129086 188956 129142
rect 189004 129086 189060 129142
rect 188796 128982 188852 129038
rect 188900 128982 188956 129038
rect 189004 128982 189060 129038
rect 188796 128878 188852 128934
rect 188900 128878 188956 128934
rect 189004 128878 189060 128934
rect 158736 99110 158792 99166
rect 158840 99110 158896 99166
rect 158944 99110 159000 99166
rect 158736 99006 158792 99062
rect 158840 99006 158896 99062
rect 158944 99006 159000 99062
rect 158736 98902 158792 98958
rect 158840 98902 158896 98958
rect 158944 98902 159000 98958
rect 184022 99110 184078 99166
rect 184022 99006 184078 99062
rect 184022 98902 184078 98958
rect 185962 99110 186018 99166
rect 186066 99110 186122 99166
rect 186170 99110 186226 99166
rect 185962 99006 186018 99062
rect 186066 99006 186122 99062
rect 186170 99006 186226 99062
rect 185962 98902 186018 98958
rect 186066 98902 186122 98958
rect 186170 98902 186226 98958
rect 184458 98450 184514 98506
rect 184458 98346 184514 98402
rect 184458 98242 184514 98298
rect 185302 98450 185358 98506
rect 185406 98450 185462 98506
rect 185510 98450 185566 98506
rect 185302 98346 185358 98402
rect 185406 98346 185462 98402
rect 185510 98346 185566 98402
rect 185302 98242 185358 98298
rect 185406 98242 185462 98298
rect 185510 98242 185566 98298
rect 188796 98450 188852 98506
rect 188900 98450 188956 98506
rect 189004 98450 189060 98506
rect 188796 98346 188852 98402
rect 188900 98346 188956 98402
rect 189004 98346 189060 98402
rect 188796 98242 188852 98298
rect 188900 98242 188956 98298
rect 189004 98242 189060 98298
rect 158736 68474 158792 68530
rect 158840 68474 158896 68530
rect 158944 68474 159000 68530
rect 158736 68370 158792 68426
rect 158840 68370 158896 68426
rect 158944 68370 159000 68426
rect 158736 68266 158792 68322
rect 158840 68266 158896 68322
rect 158944 68266 159000 68322
rect 184022 68474 184078 68530
rect 184022 68370 184078 68426
rect 184022 68266 184078 68322
rect 185962 68474 186018 68530
rect 186066 68474 186122 68530
rect 186170 68474 186226 68530
rect 185962 68370 186018 68426
rect 186066 68370 186122 68426
rect 186170 68370 186226 68426
rect 185962 68266 186018 68322
rect 186066 68266 186122 68322
rect 186170 68266 186226 68322
rect 184458 67814 184514 67870
rect 184458 67710 184514 67766
rect 184458 67606 184514 67662
rect 185302 67814 185358 67870
rect 185406 67814 185462 67870
rect 185510 67814 185566 67870
rect 185302 67710 185358 67766
rect 185406 67710 185462 67766
rect 185510 67710 185566 67766
rect 185302 67606 185358 67662
rect 185406 67606 185462 67662
rect 185510 67606 185566 67662
rect 188796 67814 188852 67870
rect 188900 67814 188956 67870
rect 189004 67814 189060 67870
rect 188796 67710 188852 67766
rect 188900 67710 188956 67766
rect 189004 67710 189060 67766
rect 188796 67606 188852 67662
rect 188900 67606 188956 67662
rect 189004 67606 189060 67662
rect 158736 37838 158792 37894
rect 158840 37838 158896 37894
rect 158944 37838 159000 37894
rect 158736 37734 158792 37790
rect 158840 37734 158896 37790
rect 158944 37734 159000 37790
rect 158736 37630 158792 37686
rect 158840 37630 158896 37686
rect 158944 37630 159000 37686
rect 161250 37838 161306 37894
rect 161250 37734 161306 37790
rect 161250 37630 161306 37686
rect 185962 37838 186018 37894
rect 186066 37838 186122 37894
rect 186170 37838 186226 37894
rect 185962 37734 186018 37790
rect 186066 37734 186122 37790
rect 186170 37734 186226 37790
rect 185962 37630 186018 37686
rect 186066 37630 186122 37686
rect 186170 37630 186226 37686
rect 185302 37178 185358 37234
rect 185406 37178 185462 37234
rect 185510 37178 185566 37234
rect 185302 37074 185358 37130
rect 185406 37074 185462 37130
rect 185510 37074 185566 37130
rect 185302 36970 185358 37026
rect 185406 36970 185462 37026
rect 185510 36970 185566 37026
rect 188796 37178 188852 37234
rect 188900 37178 188956 37234
rect 189004 37178 189060 37234
rect 188796 37074 188852 37130
rect 188900 37074 188956 37130
rect 189004 37074 189060 37130
rect 188796 36970 188852 37026
rect 188900 36970 188956 37026
rect 189004 36970 189060 37026
rect 158736 7202 158792 7258
rect 158840 7202 158896 7258
rect 158944 7202 159000 7258
rect 158736 7098 158792 7154
rect 158840 7098 158896 7154
rect 158944 7098 159000 7154
rect 158736 6994 158792 7050
rect 158840 6994 158896 7050
rect 158944 6994 159000 7050
rect 188796 6542 188852 6598
rect 188900 6542 188956 6598
rect 189004 6542 189060 6598
rect 188796 6438 188852 6494
rect 188900 6438 188956 6494
rect 189004 6438 189060 6494
rect 188796 6334 188852 6390
rect 188900 6334 188956 6390
rect 189004 6334 189060 6390
rect 189456 129746 189512 129802
rect 189560 129746 189616 129802
rect 189664 129746 189720 129802
rect 189456 129642 189512 129698
rect 189560 129642 189616 129698
rect 189664 129642 189720 129698
rect 189456 129538 189512 129594
rect 189560 129538 189616 129594
rect 189664 129538 189720 129594
rect 189456 99110 189512 99166
rect 189560 99110 189616 99166
rect 189664 99110 189720 99166
rect 189456 99006 189512 99062
rect 189560 99006 189616 99062
rect 189664 99006 189720 99062
rect 189456 98902 189512 98958
rect 189560 98902 189616 98958
rect 189664 98902 189720 98958
rect 189456 68474 189512 68530
rect 189560 68474 189616 68530
rect 189664 68474 189720 68530
rect 189456 68370 189512 68426
rect 189560 68370 189616 68426
rect 189664 68370 189720 68426
rect 189456 68266 189512 68322
rect 189560 68266 189616 68322
rect 189664 68266 189720 68322
rect 189456 37838 189512 37894
rect 189560 37838 189616 37894
rect 189664 37838 189720 37894
rect 189456 37734 189512 37790
rect 189560 37734 189616 37790
rect 189664 37734 189720 37790
rect 189456 37660 189512 37686
rect 189456 37630 189512 37660
rect 189560 37660 189616 37686
rect 189560 37630 189616 37660
rect 189664 37660 189720 37686
rect 189664 37630 189720 37660
rect 189456 7202 189512 7258
rect 189560 7202 189616 7258
rect 189664 7202 189720 7258
rect 189456 7098 189512 7154
rect 189560 7098 189616 7154
rect 189664 7098 189720 7154
rect 189456 6994 189512 7050
rect 189560 6994 189616 7050
rect 189664 6994 189720 7050
<< metal5 >>
rect 1284 129802 204796 129830
rect 1284 129746 5136 129802
rect 5192 129746 5240 129802
rect 5296 129746 5344 129802
rect 5400 129746 20038 129802
rect 20094 129746 20142 129802
rect 20198 129746 20246 129802
rect 20302 129746 35856 129802
rect 35912 129746 35960 129802
rect 36016 129746 36064 129802
rect 36120 129746 48528 129802
rect 48584 129746 49962 129802
rect 50018 129746 51414 129802
rect 51470 129746 54666 129802
rect 54722 129746 65732 129802
rect 65788 129746 66576 129802
rect 66632 129746 66680 129802
rect 66736 129746 66784 129802
rect 66840 129746 97296 129802
rect 97352 129746 97400 129802
rect 97456 129746 97504 129802
rect 97560 129746 128016 129802
rect 128072 129746 128120 129802
rect 128176 129746 128224 129802
rect 128280 129746 158736 129802
rect 158792 129746 158840 129802
rect 158896 129746 158944 129802
rect 159000 129746 184022 129802
rect 184078 129746 185962 129802
rect 186018 129746 186066 129802
rect 186122 129746 186170 129802
rect 186226 129746 189456 129802
rect 189512 129746 189560 129802
rect 189616 129746 189664 129802
rect 189720 129746 204796 129802
rect 1284 129698 204796 129746
rect 1284 129642 5136 129698
rect 5192 129642 5240 129698
rect 5296 129642 5344 129698
rect 5400 129642 20038 129698
rect 20094 129642 20142 129698
rect 20198 129642 20246 129698
rect 20302 129642 35856 129698
rect 35912 129642 35960 129698
rect 36016 129642 36064 129698
rect 36120 129642 48528 129698
rect 48584 129642 49962 129698
rect 50018 129642 51414 129698
rect 51470 129642 54666 129698
rect 54722 129642 65732 129698
rect 65788 129642 66576 129698
rect 66632 129642 66680 129698
rect 66736 129642 66784 129698
rect 66840 129642 97296 129698
rect 97352 129642 97400 129698
rect 97456 129642 97504 129698
rect 97560 129642 128016 129698
rect 128072 129642 128120 129698
rect 128176 129642 128224 129698
rect 128280 129642 158736 129698
rect 158792 129642 158840 129698
rect 158896 129642 158944 129698
rect 159000 129642 184022 129698
rect 184078 129642 185962 129698
rect 186018 129642 186066 129698
rect 186122 129642 186170 129698
rect 186226 129642 189456 129698
rect 189512 129642 189560 129698
rect 189616 129642 189664 129698
rect 189720 129642 204796 129698
rect 1284 129594 204796 129642
rect 1284 129538 5136 129594
rect 5192 129538 5240 129594
rect 5296 129538 5344 129594
rect 5400 129538 20038 129594
rect 20094 129538 20142 129594
rect 20198 129538 20246 129594
rect 20302 129538 35856 129594
rect 35912 129538 35960 129594
rect 36016 129538 36064 129594
rect 36120 129538 48528 129594
rect 48584 129538 49962 129594
rect 50018 129538 51414 129594
rect 51470 129538 54666 129594
rect 54722 129538 65732 129594
rect 65788 129538 66576 129594
rect 66632 129538 66680 129594
rect 66736 129538 66784 129594
rect 66840 129538 97296 129594
rect 97352 129538 97400 129594
rect 97456 129538 97504 129594
rect 97560 129538 128016 129594
rect 128072 129538 128120 129594
rect 128176 129538 128224 129594
rect 128280 129538 158736 129594
rect 158792 129538 158840 129594
rect 158896 129538 158944 129594
rect 159000 129538 184022 129594
rect 184078 129538 185962 129594
rect 186018 129538 186066 129594
rect 186122 129538 186170 129594
rect 186226 129538 189456 129594
rect 189512 129538 189560 129594
rect 189616 129538 189664 129594
rect 189720 129538 204796 129594
rect 1284 129510 204796 129538
rect 1284 129142 204796 129170
rect 1284 129086 4476 129142
rect 4532 129086 4580 129142
rect 4636 129086 4684 129142
rect 4740 129086 20698 129142
rect 20754 129086 20802 129142
rect 20858 129086 20906 129142
rect 20962 129086 35196 129142
rect 35252 129086 35300 129142
rect 35356 129086 35404 129142
rect 35460 129086 49598 129142
rect 49654 129086 50598 129142
rect 50654 129086 52039 129142
rect 52095 129086 60826 129142
rect 60882 129086 65296 129142
rect 65352 129086 96636 129142
rect 96692 129086 96740 129142
rect 96796 129086 96844 129142
rect 96900 129086 127356 129142
rect 127412 129086 127460 129142
rect 127516 129086 127564 129142
rect 127620 129086 158076 129142
rect 158132 129086 158180 129142
rect 158236 129086 158284 129142
rect 158340 129086 184458 129142
rect 184514 129086 185302 129142
rect 185358 129086 185406 129142
rect 185462 129086 185510 129142
rect 185566 129086 188796 129142
rect 188852 129086 188900 129142
rect 188956 129086 189004 129142
rect 189060 129086 204796 129142
rect 1284 129038 204796 129086
rect 1284 128982 4476 129038
rect 4532 128982 4580 129038
rect 4636 128982 4684 129038
rect 4740 128982 20698 129038
rect 20754 128982 20802 129038
rect 20858 128982 20906 129038
rect 20962 128982 35196 129038
rect 35252 128982 35300 129038
rect 35356 128982 35404 129038
rect 35460 128982 49598 129038
rect 49654 128982 50598 129038
rect 50654 128982 52039 129038
rect 52095 128982 60826 129038
rect 60882 128982 65296 129038
rect 65352 128982 96636 129038
rect 96692 128982 96740 129038
rect 96796 128982 96844 129038
rect 96900 128982 127356 129038
rect 127412 128982 127460 129038
rect 127516 128982 127564 129038
rect 127620 128982 158076 129038
rect 158132 128982 158180 129038
rect 158236 128982 158284 129038
rect 158340 128982 184458 129038
rect 184514 128982 185302 129038
rect 185358 128982 185406 129038
rect 185462 128982 185510 129038
rect 185566 128982 188796 129038
rect 188852 128982 188900 129038
rect 188956 128982 189004 129038
rect 189060 128982 204796 129038
rect 1284 128934 204796 128982
rect 1284 128878 4476 128934
rect 4532 128878 4580 128934
rect 4636 128878 4684 128934
rect 4740 128878 20698 128934
rect 20754 128878 20802 128934
rect 20858 128878 20906 128934
rect 20962 128878 35196 128934
rect 35252 128878 35300 128934
rect 35356 128878 35404 128934
rect 35460 128878 49598 128934
rect 49654 128878 50598 128934
rect 50654 128878 52039 128934
rect 52095 128878 60826 128934
rect 60882 128878 65296 128934
rect 65352 128878 96636 128934
rect 96692 128878 96740 128934
rect 96796 128878 96844 128934
rect 96900 128878 127356 128934
rect 127412 128878 127460 128934
rect 127516 128878 127564 128934
rect 127620 128878 158076 128934
rect 158132 128878 158180 128934
rect 158236 128878 158284 128934
rect 158340 128878 184458 128934
rect 184514 128878 185302 128934
rect 185358 128878 185406 128934
rect 185462 128878 185510 128934
rect 185566 128878 188796 128934
rect 188852 128878 188900 128934
rect 188956 128878 189004 128934
rect 189060 128878 204796 128934
rect 1284 128850 204796 128878
rect 1284 99166 204796 99194
rect 1284 99110 5136 99166
rect 5192 99110 5240 99166
rect 5296 99110 5344 99166
rect 5400 99110 20038 99166
rect 20094 99110 20142 99166
rect 20198 99110 20246 99166
rect 20302 99110 35856 99166
rect 35912 99110 35960 99166
rect 36016 99110 36064 99166
rect 36120 99110 48528 99166
rect 48584 99110 49962 99166
rect 50018 99110 51414 99166
rect 51470 99110 54666 99166
rect 54722 99110 65732 99166
rect 65788 99110 66576 99166
rect 66632 99110 66680 99166
rect 66736 99110 66784 99166
rect 66840 99110 97296 99166
rect 97352 99110 97400 99166
rect 97456 99110 97504 99166
rect 97560 99110 128016 99166
rect 128072 99110 128120 99166
rect 128176 99110 128224 99166
rect 128280 99110 158736 99166
rect 158792 99110 158840 99166
rect 158896 99110 158944 99166
rect 159000 99110 184022 99166
rect 184078 99110 185962 99166
rect 186018 99110 186066 99166
rect 186122 99110 186170 99166
rect 186226 99110 189456 99166
rect 189512 99110 189560 99166
rect 189616 99110 189664 99166
rect 189720 99110 204796 99166
rect 1284 99062 204796 99110
rect 1284 99006 5136 99062
rect 5192 99006 5240 99062
rect 5296 99006 5344 99062
rect 5400 99006 20038 99062
rect 20094 99006 20142 99062
rect 20198 99006 20246 99062
rect 20302 99006 35856 99062
rect 35912 99006 35960 99062
rect 36016 99006 36064 99062
rect 36120 99006 48528 99062
rect 48584 99006 49962 99062
rect 50018 99006 51414 99062
rect 51470 99006 54666 99062
rect 54722 99006 65732 99062
rect 65788 99006 66576 99062
rect 66632 99006 66680 99062
rect 66736 99006 66784 99062
rect 66840 99006 97296 99062
rect 97352 99006 97400 99062
rect 97456 99006 97504 99062
rect 97560 99006 128016 99062
rect 128072 99006 128120 99062
rect 128176 99006 128224 99062
rect 128280 99006 158736 99062
rect 158792 99006 158840 99062
rect 158896 99006 158944 99062
rect 159000 99006 184022 99062
rect 184078 99006 185962 99062
rect 186018 99006 186066 99062
rect 186122 99006 186170 99062
rect 186226 99006 189456 99062
rect 189512 99006 189560 99062
rect 189616 99006 189664 99062
rect 189720 99006 204796 99062
rect 1284 98958 204796 99006
rect 1284 98902 5136 98958
rect 5192 98902 5240 98958
rect 5296 98902 5344 98958
rect 5400 98902 20038 98958
rect 20094 98902 20142 98958
rect 20198 98902 20246 98958
rect 20302 98902 35856 98958
rect 35912 98902 35960 98958
rect 36016 98902 36064 98958
rect 36120 98902 48528 98958
rect 48584 98902 49962 98958
rect 50018 98902 51414 98958
rect 51470 98902 54666 98958
rect 54722 98902 65732 98958
rect 65788 98902 66576 98958
rect 66632 98902 66680 98958
rect 66736 98902 66784 98958
rect 66840 98902 97296 98958
rect 97352 98902 97400 98958
rect 97456 98902 97504 98958
rect 97560 98902 128016 98958
rect 128072 98902 128120 98958
rect 128176 98902 128224 98958
rect 128280 98902 158736 98958
rect 158792 98902 158840 98958
rect 158896 98902 158944 98958
rect 159000 98902 184022 98958
rect 184078 98902 185962 98958
rect 186018 98902 186066 98958
rect 186122 98902 186170 98958
rect 186226 98902 189456 98958
rect 189512 98902 189560 98958
rect 189616 98902 189664 98958
rect 189720 98902 204796 98958
rect 1284 98874 204796 98902
rect 1284 98506 204796 98534
rect 1284 98450 4476 98506
rect 4532 98450 4580 98506
rect 4636 98450 4684 98506
rect 4740 98450 20698 98506
rect 20754 98450 20802 98506
rect 20858 98450 20906 98506
rect 20962 98450 35196 98506
rect 35252 98450 35300 98506
rect 35356 98450 35404 98506
rect 35460 98450 49598 98506
rect 49654 98450 50598 98506
rect 50654 98450 52039 98506
rect 52095 98450 60826 98506
rect 60882 98450 65296 98506
rect 65352 98450 96636 98506
rect 96692 98450 96740 98506
rect 96796 98450 96844 98506
rect 96900 98450 127356 98506
rect 127412 98450 127460 98506
rect 127516 98450 127564 98506
rect 127620 98450 158076 98506
rect 158132 98450 158180 98506
rect 158236 98450 158284 98506
rect 158340 98450 184458 98506
rect 184514 98450 185302 98506
rect 185358 98450 185406 98506
rect 185462 98450 185510 98506
rect 185566 98450 188796 98506
rect 188852 98450 188900 98506
rect 188956 98450 189004 98506
rect 189060 98450 204796 98506
rect 1284 98402 204796 98450
rect 1284 98346 4476 98402
rect 4532 98346 4580 98402
rect 4636 98346 4684 98402
rect 4740 98346 20698 98402
rect 20754 98346 20802 98402
rect 20858 98346 20906 98402
rect 20962 98346 35196 98402
rect 35252 98346 35300 98402
rect 35356 98346 35404 98402
rect 35460 98346 49598 98402
rect 49654 98346 50598 98402
rect 50654 98346 52039 98402
rect 52095 98346 60826 98402
rect 60882 98346 65296 98402
rect 65352 98346 96636 98402
rect 96692 98346 96740 98402
rect 96796 98346 96844 98402
rect 96900 98346 127356 98402
rect 127412 98346 127460 98402
rect 127516 98346 127564 98402
rect 127620 98346 158076 98402
rect 158132 98346 158180 98402
rect 158236 98346 158284 98402
rect 158340 98346 184458 98402
rect 184514 98346 185302 98402
rect 185358 98346 185406 98402
rect 185462 98346 185510 98402
rect 185566 98346 188796 98402
rect 188852 98346 188900 98402
rect 188956 98346 189004 98402
rect 189060 98346 204796 98402
rect 1284 98298 204796 98346
rect 1284 98242 4476 98298
rect 4532 98242 4580 98298
rect 4636 98242 4684 98298
rect 4740 98242 20698 98298
rect 20754 98242 20802 98298
rect 20858 98242 20906 98298
rect 20962 98242 35196 98298
rect 35252 98242 35300 98298
rect 35356 98242 35404 98298
rect 35460 98242 49598 98298
rect 49654 98242 50598 98298
rect 50654 98242 52039 98298
rect 52095 98242 60826 98298
rect 60882 98242 65296 98298
rect 65352 98242 96636 98298
rect 96692 98242 96740 98298
rect 96796 98242 96844 98298
rect 96900 98242 127356 98298
rect 127412 98242 127460 98298
rect 127516 98242 127564 98298
rect 127620 98242 158076 98298
rect 158132 98242 158180 98298
rect 158236 98242 158284 98298
rect 158340 98242 184458 98298
rect 184514 98242 185302 98298
rect 185358 98242 185406 98298
rect 185462 98242 185510 98298
rect 185566 98242 188796 98298
rect 188852 98242 188900 98298
rect 188956 98242 189004 98298
rect 189060 98242 204796 98298
rect 1284 98214 204796 98242
rect 1284 68530 204796 68558
rect 1284 68474 5136 68530
rect 5192 68474 5240 68530
rect 5296 68474 5344 68530
rect 5400 68474 20038 68530
rect 20094 68474 20142 68530
rect 20198 68474 20246 68530
rect 20302 68474 35856 68530
rect 35912 68474 35960 68530
rect 36016 68474 36064 68530
rect 36120 68474 48528 68530
rect 48584 68474 49962 68530
rect 50018 68474 51414 68530
rect 51470 68474 54666 68530
rect 54722 68474 65732 68530
rect 65788 68474 66576 68530
rect 66632 68474 66680 68530
rect 66736 68474 66784 68530
rect 66840 68474 97296 68530
rect 97352 68474 97400 68530
rect 97456 68474 97504 68530
rect 97560 68474 128016 68530
rect 128072 68474 128120 68530
rect 128176 68474 128224 68530
rect 128280 68474 158736 68530
rect 158792 68474 158840 68530
rect 158896 68474 158944 68530
rect 159000 68474 184022 68530
rect 184078 68474 185962 68530
rect 186018 68474 186066 68530
rect 186122 68474 186170 68530
rect 186226 68474 189456 68530
rect 189512 68474 189560 68530
rect 189616 68474 189664 68530
rect 189720 68474 204796 68530
rect 1284 68459 204796 68474
rect 1284 68426 44562 68459
rect 1284 68370 5136 68426
rect 5192 68370 5240 68426
rect 5296 68370 5344 68426
rect 5400 68370 20038 68426
rect 20094 68370 20142 68426
rect 20198 68370 20246 68426
rect 20302 68370 35856 68426
rect 35912 68370 35960 68426
rect 36016 68370 36064 68426
rect 36120 68403 44562 68426
rect 44618 68426 204796 68459
rect 44618 68403 48528 68426
rect 36120 68370 48528 68403
rect 48584 68370 49962 68426
rect 50018 68370 51414 68426
rect 51470 68370 54666 68426
rect 54722 68370 65732 68426
rect 65788 68370 66576 68426
rect 66632 68370 66680 68426
rect 66736 68370 66784 68426
rect 66840 68370 97296 68426
rect 97352 68370 97400 68426
rect 97456 68370 97504 68426
rect 97560 68370 128016 68426
rect 128072 68370 128120 68426
rect 128176 68370 128224 68426
rect 128280 68370 158736 68426
rect 158792 68370 158840 68426
rect 158896 68370 158944 68426
rect 159000 68370 184022 68426
rect 184078 68370 185962 68426
rect 186018 68370 186066 68426
rect 186122 68370 186170 68426
rect 186226 68370 189456 68426
rect 189512 68370 189560 68426
rect 189616 68370 189664 68426
rect 189720 68370 204796 68426
rect 1284 68355 204796 68370
rect 1284 68341 44562 68355
rect 1284 68322 42582 68341
rect 1284 68266 5136 68322
rect 5192 68266 5240 68322
rect 5296 68266 5344 68322
rect 5400 68266 20038 68322
rect 20094 68266 20142 68322
rect 20198 68266 20246 68322
rect 20302 68266 35856 68322
rect 35912 68266 35960 68322
rect 36016 68266 36064 68322
rect 36120 68285 42582 68322
rect 42638 68299 44562 68341
rect 44618 68322 204796 68355
rect 44618 68299 48528 68322
rect 42638 68285 48528 68299
rect 36120 68266 48528 68285
rect 48584 68266 49962 68322
rect 50018 68266 51414 68322
rect 51470 68266 54666 68322
rect 54722 68266 65732 68322
rect 65788 68266 66576 68322
rect 66632 68266 66680 68322
rect 66736 68266 66784 68322
rect 66840 68266 97296 68322
rect 97352 68266 97400 68322
rect 97456 68266 97504 68322
rect 97560 68266 128016 68322
rect 128072 68266 128120 68322
rect 128176 68266 128224 68322
rect 128280 68266 158736 68322
rect 158792 68266 158840 68322
rect 158896 68266 158944 68322
rect 159000 68266 184022 68322
rect 184078 68266 185962 68322
rect 186018 68266 186066 68322
rect 186122 68266 186170 68322
rect 186226 68266 189456 68322
rect 189512 68266 189560 68322
rect 189616 68266 189664 68322
rect 189720 68266 204796 68322
rect 1284 68238 204796 68266
rect 1284 67870 204796 67898
rect 1284 67814 4476 67870
rect 4532 67814 4580 67870
rect 4636 67814 4684 67870
rect 4740 67814 20698 67870
rect 20754 67814 20802 67870
rect 20858 67814 20906 67870
rect 20962 67814 35196 67870
rect 35252 67814 35300 67870
rect 35356 67814 35404 67870
rect 35460 67855 49598 67870
rect 35460 67814 44694 67855
rect 1284 67799 44694 67814
rect 44750 67799 46014 67855
rect 46070 67814 49598 67855
rect 49654 67814 50598 67870
rect 50654 67814 52039 67870
rect 52095 67814 60826 67870
rect 60882 67814 65296 67870
rect 65352 67814 96636 67870
rect 96692 67814 96740 67870
rect 96796 67814 96844 67870
rect 96900 67814 127356 67870
rect 127412 67814 127460 67870
rect 127516 67814 127564 67870
rect 127620 67814 158076 67870
rect 158132 67814 158180 67870
rect 158236 67814 158284 67870
rect 158340 67814 184458 67870
rect 184514 67814 185302 67870
rect 185358 67814 185406 67870
rect 185462 67814 185510 67870
rect 185566 67814 188796 67870
rect 188852 67814 188900 67870
rect 188956 67814 189004 67870
rect 189060 67814 204796 67870
rect 46070 67799 204796 67814
rect 1284 67766 204796 67799
rect 1284 67710 4476 67766
rect 4532 67710 4580 67766
rect 4636 67710 4684 67766
rect 4740 67710 20698 67766
rect 20754 67710 20802 67766
rect 20858 67710 20906 67766
rect 20962 67710 35196 67766
rect 35252 67710 35300 67766
rect 35356 67710 35404 67766
rect 35460 67751 49598 67766
rect 35460 67710 44694 67751
rect 1284 67695 44694 67710
rect 44750 67695 46014 67751
rect 46070 67710 49598 67751
rect 49654 67710 50598 67766
rect 50654 67710 52039 67766
rect 52095 67710 60826 67766
rect 60882 67710 65296 67766
rect 65352 67710 96636 67766
rect 96692 67710 96740 67766
rect 96796 67710 96844 67766
rect 96900 67710 127356 67766
rect 127412 67710 127460 67766
rect 127516 67710 127564 67766
rect 127620 67710 158076 67766
rect 158132 67710 158180 67766
rect 158236 67710 158284 67766
rect 158340 67710 184458 67766
rect 184514 67710 185302 67766
rect 185358 67710 185406 67766
rect 185462 67710 185510 67766
rect 185566 67710 188796 67766
rect 188852 67710 188900 67766
rect 188956 67710 189004 67766
rect 189060 67710 204796 67766
rect 46070 67695 204796 67710
rect 1284 67662 204796 67695
rect 1284 67606 4476 67662
rect 4532 67606 4580 67662
rect 4636 67606 4684 67662
rect 4740 67606 20698 67662
rect 20754 67606 20802 67662
rect 20858 67606 20906 67662
rect 20962 67606 35196 67662
rect 35252 67606 35300 67662
rect 35356 67606 35404 67662
rect 35460 67606 49598 67662
rect 49654 67606 50598 67662
rect 50654 67606 52039 67662
rect 52095 67606 60826 67662
rect 60882 67606 65296 67662
rect 65352 67606 96636 67662
rect 96692 67606 96740 67662
rect 96796 67606 96844 67662
rect 96900 67606 127356 67662
rect 127412 67606 127460 67662
rect 127516 67606 127564 67662
rect 127620 67606 158076 67662
rect 158132 67606 158180 67662
rect 158236 67606 158284 67662
rect 158340 67606 184458 67662
rect 184514 67606 185302 67662
rect 185358 67606 185406 67662
rect 185462 67606 185510 67662
rect 185566 67606 188796 67662
rect 188852 67606 188900 67662
rect 188956 67606 189004 67662
rect 189060 67606 204796 67662
rect 1284 67578 204796 67606
rect 1284 37894 204796 37922
rect 1284 37838 5136 37894
rect 5192 37838 5240 37894
rect 5296 37838 5344 37894
rect 5400 37838 20038 37894
rect 20094 37838 20142 37894
rect 20198 37838 20246 37894
rect 20302 37838 29062 37894
rect 29118 37838 35856 37894
rect 35912 37838 35960 37894
rect 36016 37838 36064 37894
rect 36120 37838 43728 37894
rect 43784 37838 45970 37894
rect 46026 37838 47652 37894
rect 47708 37838 66576 37894
rect 66632 37838 66680 37894
rect 66736 37838 66784 37894
rect 66840 37838 97296 37894
rect 97352 37838 97400 37894
rect 97456 37838 97504 37894
rect 97560 37838 128016 37894
rect 128072 37838 128120 37894
rect 128176 37838 128224 37894
rect 128280 37838 158736 37894
rect 158792 37838 158840 37894
rect 158896 37838 158944 37894
rect 159000 37838 161250 37894
rect 161306 37838 185962 37894
rect 186018 37838 186066 37894
rect 186122 37838 186170 37894
rect 186226 37838 189456 37894
rect 189512 37838 189560 37894
rect 189616 37838 189664 37894
rect 189720 37838 204796 37894
rect 1284 37790 204796 37838
rect 1284 37734 5136 37790
rect 5192 37734 5240 37790
rect 5296 37734 5344 37790
rect 5400 37734 20038 37790
rect 20094 37734 20142 37790
rect 20198 37734 20246 37790
rect 20302 37734 29062 37790
rect 29118 37734 35856 37790
rect 35912 37734 35960 37790
rect 36016 37734 36064 37790
rect 36120 37734 43728 37790
rect 43784 37734 45970 37790
rect 46026 37734 47652 37790
rect 47708 37734 66576 37790
rect 66632 37734 66680 37790
rect 66736 37734 66784 37790
rect 66840 37734 97296 37790
rect 97352 37734 97400 37790
rect 97456 37734 97504 37790
rect 97560 37734 128016 37790
rect 128072 37734 128120 37790
rect 128176 37734 128224 37790
rect 128280 37734 158736 37790
rect 158792 37734 158840 37790
rect 158896 37734 158944 37790
rect 159000 37734 161250 37790
rect 161306 37734 185962 37790
rect 186018 37734 186066 37790
rect 186122 37734 186170 37790
rect 186226 37734 189456 37790
rect 189512 37734 189560 37790
rect 189616 37734 189664 37790
rect 189720 37734 204796 37790
rect 1284 37686 204796 37734
rect 1284 37630 5136 37686
rect 5192 37630 5240 37686
rect 5296 37630 5344 37686
rect 5400 37630 20038 37686
rect 20094 37630 20142 37686
rect 20198 37630 20246 37686
rect 20302 37630 29062 37686
rect 29118 37630 35856 37686
rect 35912 37630 35960 37686
rect 36016 37630 36064 37686
rect 36120 37630 43728 37686
rect 43784 37630 45970 37686
rect 46026 37630 47652 37686
rect 47708 37630 66576 37686
rect 66632 37630 66680 37686
rect 66736 37630 66784 37686
rect 66840 37630 97296 37686
rect 97352 37630 97400 37686
rect 97456 37630 97504 37686
rect 97560 37630 128016 37686
rect 128072 37630 128120 37686
rect 128176 37630 128224 37686
rect 128280 37630 158736 37686
rect 158792 37630 158840 37686
rect 158896 37630 158944 37686
rect 159000 37630 161250 37686
rect 161306 37630 185962 37686
rect 186018 37630 186066 37686
rect 186122 37630 186170 37686
rect 186226 37630 189456 37686
rect 189512 37630 189560 37686
rect 189616 37630 189664 37686
rect 189720 37630 204796 37686
rect 1284 37602 204796 37630
rect 1284 37234 204796 37262
rect 1284 37178 4476 37234
rect 4532 37178 4580 37234
rect 4636 37178 4684 37234
rect 4740 37178 20698 37234
rect 20754 37178 20802 37234
rect 20858 37178 20906 37234
rect 20962 37178 35196 37234
rect 35252 37178 35300 37234
rect 35356 37178 35404 37234
rect 35460 37178 40074 37234
rect 40130 37178 44384 37234
rect 44440 37178 47294 37234
rect 47350 37178 48308 37234
rect 48364 37178 127356 37234
rect 127412 37178 127460 37234
rect 127516 37178 127564 37234
rect 127620 37178 130890 37234
rect 130946 37178 158076 37234
rect 158132 37178 158180 37234
rect 158236 37178 158284 37234
rect 158340 37178 185302 37234
rect 185358 37178 185406 37234
rect 185462 37178 185510 37234
rect 185566 37178 188796 37234
rect 188852 37178 188900 37234
rect 188956 37178 189004 37234
rect 189060 37178 204796 37234
rect 1284 37130 204796 37178
rect 1284 37074 4476 37130
rect 4532 37074 4580 37130
rect 4636 37074 4684 37130
rect 4740 37074 20698 37130
rect 20754 37074 20802 37130
rect 20858 37074 20906 37130
rect 20962 37074 35196 37130
rect 35252 37074 35300 37130
rect 35356 37074 35404 37130
rect 35460 37074 40074 37130
rect 40130 37074 44384 37130
rect 44440 37074 47294 37130
rect 47350 37074 48308 37130
rect 48364 37074 127356 37130
rect 127412 37074 127460 37130
rect 127516 37074 127564 37130
rect 127620 37074 130890 37130
rect 130946 37074 158076 37130
rect 158132 37074 158180 37130
rect 158236 37074 158284 37130
rect 158340 37074 185302 37130
rect 185358 37074 185406 37130
rect 185462 37074 185510 37130
rect 185566 37074 188796 37130
rect 188852 37074 188900 37130
rect 188956 37074 189004 37130
rect 189060 37074 204796 37130
rect 1284 37026 204796 37074
rect 1284 36970 4476 37026
rect 4532 36970 4580 37026
rect 4636 36970 4684 37026
rect 4740 36970 20698 37026
rect 20754 36970 20802 37026
rect 20858 36970 20906 37026
rect 20962 36970 35196 37026
rect 35252 36970 35300 37026
rect 35356 36970 35404 37026
rect 35460 36970 40074 37026
rect 40130 36970 44384 37026
rect 44440 36970 47294 37026
rect 47350 36970 48308 37026
rect 48364 36970 127356 37026
rect 127412 36970 127460 37026
rect 127516 36970 127564 37026
rect 127620 36970 130890 37026
rect 130946 36970 158076 37026
rect 158132 36970 158180 37026
rect 158236 36970 158284 37026
rect 158340 36970 185302 37026
rect 185358 36970 185406 37026
rect 185462 36970 185510 37026
rect 185566 36970 188796 37026
rect 188852 36970 188900 37026
rect 188956 36970 189004 37026
rect 189060 36970 204796 37026
rect 1284 36942 204796 36970
rect 1284 7258 204796 7286
rect 1284 7202 5136 7258
rect 5192 7202 5240 7258
rect 5296 7202 5344 7258
rect 5400 7202 35856 7258
rect 35912 7202 35960 7258
rect 36016 7202 36064 7258
rect 36120 7202 66576 7258
rect 66632 7202 66680 7258
rect 66736 7202 66784 7258
rect 66840 7202 97296 7258
rect 97352 7202 97400 7258
rect 97456 7202 97504 7258
rect 97560 7202 128016 7258
rect 128072 7202 128120 7258
rect 128176 7202 128224 7258
rect 128280 7202 158736 7258
rect 158792 7202 158840 7258
rect 158896 7202 158944 7258
rect 159000 7202 189456 7258
rect 189512 7202 189560 7258
rect 189616 7202 189664 7258
rect 189720 7202 204796 7258
rect 1284 7154 204796 7202
rect 1284 7098 5136 7154
rect 5192 7098 5240 7154
rect 5296 7098 5344 7154
rect 5400 7098 35856 7154
rect 35912 7098 35960 7154
rect 36016 7098 36064 7154
rect 36120 7098 66576 7154
rect 66632 7098 66680 7154
rect 66736 7098 66784 7154
rect 66840 7098 97296 7154
rect 97352 7098 97400 7154
rect 97456 7098 97504 7154
rect 97560 7098 128016 7154
rect 128072 7098 128120 7154
rect 128176 7098 128224 7154
rect 128280 7098 158736 7154
rect 158792 7098 158840 7154
rect 158896 7098 158944 7154
rect 159000 7098 189456 7154
rect 189512 7098 189560 7154
rect 189616 7098 189664 7154
rect 189720 7098 204796 7154
rect 1284 7050 204796 7098
rect 1284 6994 5136 7050
rect 5192 6994 5240 7050
rect 5296 6994 5344 7050
rect 5400 6994 35856 7050
rect 35912 6994 35960 7050
rect 36016 6994 36064 7050
rect 36120 6994 66576 7050
rect 66632 6994 66680 7050
rect 66736 6994 66784 7050
rect 66840 6994 97296 7050
rect 97352 6994 97400 7050
rect 97456 6994 97504 7050
rect 97560 6994 128016 7050
rect 128072 6994 128120 7050
rect 128176 6994 128224 7050
rect 128280 6994 158736 7050
rect 158792 6994 158840 7050
rect 158896 6994 158944 7050
rect 159000 6994 189456 7050
rect 189512 6994 189560 7050
rect 189616 6994 189664 7050
rect 189720 6994 204796 7050
rect 1284 6966 204796 6994
rect 1284 6598 204796 6626
rect 1284 6542 4476 6598
rect 4532 6542 4580 6598
rect 4636 6542 4684 6598
rect 4740 6542 35196 6598
rect 35252 6542 35300 6598
rect 35356 6542 35404 6598
rect 35460 6542 65916 6598
rect 65972 6542 66020 6598
rect 66076 6542 66124 6598
rect 66180 6542 96636 6598
rect 96692 6542 96740 6598
rect 96796 6542 96844 6598
rect 96900 6542 127356 6598
rect 127412 6542 127460 6598
rect 127516 6542 127564 6598
rect 127620 6542 158076 6598
rect 158132 6542 158180 6598
rect 158236 6542 158284 6598
rect 158340 6542 188796 6598
rect 188852 6542 188900 6598
rect 188956 6542 189004 6598
rect 189060 6542 204796 6598
rect 1284 6494 204796 6542
rect 1284 6438 4476 6494
rect 4532 6438 4580 6494
rect 4636 6438 4684 6494
rect 4740 6438 35196 6494
rect 35252 6438 35300 6494
rect 35356 6438 35404 6494
rect 35460 6438 65916 6494
rect 65972 6438 66020 6494
rect 66076 6438 66124 6494
rect 66180 6438 96636 6494
rect 96692 6438 96740 6494
rect 96796 6438 96844 6494
rect 96900 6438 127356 6494
rect 127412 6438 127460 6494
rect 127516 6438 127564 6494
rect 127620 6438 158076 6494
rect 158132 6438 158180 6494
rect 158236 6438 158284 6494
rect 158340 6438 188796 6494
rect 188852 6438 188900 6494
rect 188956 6438 189004 6494
rect 189060 6438 204796 6494
rect 1284 6390 204796 6438
rect 1284 6334 4476 6390
rect 4532 6334 4580 6390
rect 4636 6334 4684 6390
rect 4740 6334 35196 6390
rect 35252 6334 35300 6390
rect 35356 6334 35404 6390
rect 35460 6334 65916 6390
rect 65972 6334 66020 6390
rect 66076 6334 66124 6390
rect 66180 6334 96636 6390
rect 96692 6334 96740 6390
rect 96796 6334 96844 6390
rect 96900 6334 127356 6390
rect 127412 6334 127460 6390
rect 127516 6334 127564 6390
rect 127620 6334 158076 6390
rect 158132 6334 158180 6390
rect 158236 6334 158284 6390
rect 158340 6334 188796 6390
rect 188852 6334 188900 6390
rect 188956 6334 189004 6390
rect 189060 6334 204796 6390
rect 1284 6306 204796 6334
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[0] pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 44688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[1]
timestamp 1694700623
transform 1 0 48160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[2]
timestamp 1694700623
transform 1 0 51520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[3]
timestamp 1694700623
transform 1 0 55104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[4]
timestamp 1694700623
transform 1 0 17472 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[5]
timestamp 1694700623
transform 1 0 17472 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[6]
timestamp 1694700623
transform 1 0 17472 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[7]
timestamp 1694700623
transform -1 0 17696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[8]
timestamp 1694700623
transform -1 0 17696 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_addr0[9]
timestamp 1694700623
transform -1 0 17696 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_clk0
timestamp 1694700623
transform -1 0 17696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_csb0
timestamp 1694700623
transform -1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[0]
timestamp 1694700623
transform -1 0 59136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[1]
timestamp 1694700623
transform -1 0 62048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[2]
timestamp 1694700623
transform -1 0 65520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[3]
timestamp 1694700623
transform -1 0 68880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[4]
timestamp 1694700623
transform 1 0 72128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[5]
timestamp 1694700623
transform 1 0 75488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[6]
timestamp 1694700623
transform 1 0 78960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_din0[7]
timestamp 1694700623
transform 1 0 82320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[0]
timestamp 1694700623
transform 1 0 67872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[1]
timestamp 1694700623
transform -1 0 82992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[2]
timestamp 1694700623
transform -1 0 97216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[3]
timestamp 1694700623
transform -1 0 111328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[4]
timestamp 1694700623
transform -1 0 125664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[5]
timestamp 1694700623
transform -1 0 140112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[6]
timestamp 1694700623
transform -1 0 154448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_dout0[7]
timestamp 1694700623
transform 1 0 188720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_gf180_sram_8x1024_web0
timestamp 1694700623
transform -1 0 17696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1694700623
transform -1 0 110544 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1694700623
transform 1 0 89376 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1694700623
transform 1 0 66528 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1694700623
transform 1 0 43680 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1694700623
transform -1 0 19152 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1694700623
transform 1 0 1792 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1694700623
transform 1 0 1792 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1694700623
transform 1 0 1792 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1694700623
transform 1 0 1792 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1694700623
transform 1 0 1792 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1694700623
transform 1 0 2464 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1694700623
transform 1 0 2464 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1694700623
transform 1 0 2464 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1694700623
transform 1 0 2464 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1694700623
transform 1 0 1792 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1694700623
transform 1 0 1792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1694700623
transform 1 0 2464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1694700623
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1694700623
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1694700623
transform 1 0 157920 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1694700623
transform 1 0 135072 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1694700623
transform 1 0 204288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1694700623
transform 1 0 201376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1694700623
transform 1 0 203952 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output25_I
timestamp 1694700623
transform 1 0 203952 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1694700623
transform 1 0 203728 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1694700623
transform 1 0 201040 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output28_I
timestamp 1694700623
transform 1 0 197456 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output29_I
timestamp 1694700623
transform 1 0 174608 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_6 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 2016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_22 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 3808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_30 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1694700623
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1694700623
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1694700623
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1694700623
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1694700623
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1694700623
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274
timestamp 1694700623
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_290
timestamp 1694700623
transform 1 0 33824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_294 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 34272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_299
timestamp 1694700623
transform 1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1694700623
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1694700623
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1694700623
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1694700623
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1694700623
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1694700623
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_478
timestamp 1694700623
transform 1 0 54880 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_512
timestamp 1694700623
transform 1 0 58688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_546
timestamp 1694700623
transform 1 0 62496 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_580
timestamp 1694700623
transform 1 0 66304 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_614
timestamp 1694700623
transform 1 0 70112 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_648
timestamp 1694700623
transform 1 0 73920 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_682
timestamp 1694700623
transform 1 0 77728 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_716
timestamp 1694700623
transform 1 0 81536 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_750
timestamp 1694700623
transform 1 0 85344 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_784
timestamp 1694700623
transform 1 0 89152 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_818
timestamp 1694700623
transform 1 0 92960 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_852
timestamp 1694700623
transform 1 0 96768 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_886
timestamp 1694700623
transform 1 0 100576 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_902
timestamp 1694700623
transform 1 0 102368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_906
timestamp 1694700623
transform 1 0 102816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_911
timestamp 1694700623
transform 1 0 103376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_915
timestamp 1694700623
transform 1 0 103824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_917
timestamp 1694700623
transform 1 0 104048 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_920
timestamp 1694700623
transform 1 0 104384 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_954
timestamp 1694700623
transform 1 0 108192 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_988
timestamp 1694700623
transform 1 0 112000 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1022
timestamp 1694700623
transform 1 0 115808 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1056
timestamp 1694700623
transform 1 0 119616 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1090
timestamp 1694700623
transform 1 0 123424 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1124
timestamp 1694700623
transform 1 0 127232 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1158
timestamp 1694700623
transform 1 0 131040 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1192
timestamp 1694700623
transform 1 0 134848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1226
timestamp 1694700623
transform 1 0 138656 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1260
timestamp 1694700623
transform 1 0 142464 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1294
timestamp 1694700623
transform 1 0 146272 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1328
timestamp 1694700623
transform 1 0 150080 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1362
timestamp 1694700623
transform 1 0 153888 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1396
timestamp 1694700623
transform 1 0 157696 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1430
timestamp 1694700623
transform 1 0 161504 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1464
timestamp 1694700623
transform 1 0 165312 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1498
timestamp 1694700623
transform 1 0 169120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1514
timestamp 1694700623
transform 1 0 170912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1518
timestamp 1694700623
transform 1 0 171360 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1523
timestamp 1694700623
transform 1 0 171920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1527
timestamp 1694700623
transform 1 0 172368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1529
timestamp 1694700623
transform 1 0 172592 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1532
timestamp 1694700623
transform 1 0 172928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1566
timestamp 1694700623
transform 1 0 176736 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1600
timestamp 1694700623
transform 1 0 180544 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1634
timestamp 1694700623
transform 1 0 184352 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1668
timestamp 1694700623
transform 1 0 188160 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1702
timestamp 1694700623
transform 1 0 191968 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1736
timestamp 1694700623
transform 1 0 195776 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_1770
timestamp 1694700623
transform 1 0 199584 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1804
timestamp 1694700623
transform 1 0 203392 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1812
timestamp 1694700623
transform 1 0 204288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1694700623
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1694700623
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1694700623
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1694700623
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1694700623
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1694700623
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1694700623
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1694700623
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1694700623
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1694700623
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1694700623
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1694700623
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1694700623
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_492
timestamp 1694700623
transform 1 0 56448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_556
timestamp 1694700623
transform 1 0 63616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_562
timestamp 1694700623
transform 1 0 64288 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_626
timestamp 1694700623
transform 1 0 71456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_632
timestamp 1694700623
transform 1 0 72128 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_696
timestamp 1694700623
transform 1 0 79296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_702
timestamp 1694700623
transform 1 0 79968 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_766
timestamp 1694700623
transform 1 0 87136 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_772
timestamp 1694700623
transform 1 0 87808 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_836
timestamp 1694700623
transform 1 0 94976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_842
timestamp 1694700623
transform 1 0 95648 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_906
timestamp 1694700623
transform 1 0 102816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_912
timestamp 1694700623
transform 1 0 103488 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_976
timestamp 1694700623
transform 1 0 110656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_982
timestamp 1694700623
transform 1 0 111328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1046
timestamp 1694700623
transform 1 0 118496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1052
timestamp 1694700623
transform 1 0 119168 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1116
timestamp 1694700623
transform 1 0 126336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1122
timestamp 1694700623
transform 1 0 127008 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1186
timestamp 1694700623
transform 1 0 134176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1192
timestamp 1694700623
transform 1 0 134848 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1256
timestamp 1694700623
transform 1 0 142016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1262
timestamp 1694700623
transform 1 0 142688 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1326
timestamp 1694700623
transform 1 0 149856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1332
timestamp 1694700623
transform 1 0 150528 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1396
timestamp 1694700623
transform 1 0 157696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1402
timestamp 1694700623
transform 1 0 158368 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1466
timestamp 1694700623
transform 1 0 165536 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1472
timestamp 1694700623
transform 1 0 166208 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1536
timestamp 1694700623
transform 1 0 173376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1542
timestamp 1694700623
transform 1 0 174048 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1606
timestamp 1694700623
transform 1 0 181216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1612
timestamp 1694700623
transform 1 0 181888 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1676
timestamp 1694700623
transform 1 0 189056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1682
timestamp 1694700623
transform 1 0 189728 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1746
timestamp 1694700623
transform 1 0 196896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_1752
timestamp 1694700623
transform 1 0 197568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_1784
timestamp 1694700623
transform 1 0 201152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1800
timestamp 1694700623
transform 1 0 202944 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1808
timestamp 1694700623
transform 1 0 203840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1812
timestamp 1694700623
transform 1 0 204288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1694700623
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1694700623
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1694700623
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1694700623
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1694700623
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1694700623
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1694700623
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1694700623
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1694700623
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1694700623
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1694700623
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1694700623
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1694700623
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1694700623
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1694700623
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1694700623
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_527
timestamp 1694700623
transform 1 0 60368 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_591
timestamp 1694700623
transform 1 0 67536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_597
timestamp 1694700623
transform 1 0 68208 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_661
timestamp 1694700623
transform 1 0 75376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_667
timestamp 1694700623
transform 1 0 76048 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_731
timestamp 1694700623
transform 1 0 83216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_737
timestamp 1694700623
transform 1 0 83888 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_801
timestamp 1694700623
transform 1 0 91056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_807
timestamp 1694700623
transform 1 0 91728 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_871
timestamp 1694700623
transform 1 0 98896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_877
timestamp 1694700623
transform 1 0 99568 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_941
timestamp 1694700623
transform 1 0 106736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_947
timestamp 1694700623
transform 1 0 107408 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1011
timestamp 1694700623
transform 1 0 114576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1017
timestamp 1694700623
transform 1 0 115248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1081
timestamp 1694700623
transform 1 0 122416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1087
timestamp 1694700623
transform 1 0 123088 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1151
timestamp 1694700623
transform 1 0 130256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1157
timestamp 1694700623
transform 1 0 130928 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1221
timestamp 1694700623
transform 1 0 138096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1227
timestamp 1694700623
transform 1 0 138768 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1291
timestamp 1694700623
transform 1 0 145936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1297
timestamp 1694700623
transform 1 0 146608 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1361
timestamp 1694700623
transform 1 0 153776 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1367
timestamp 1694700623
transform 1 0 154448 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1431
timestamp 1694700623
transform 1 0 161616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1437
timestamp 1694700623
transform 1 0 162288 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1501
timestamp 1694700623
transform 1 0 169456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1507
timestamp 1694700623
transform 1 0 170128 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1571
timestamp 1694700623
transform 1 0 177296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1577
timestamp 1694700623
transform 1 0 177968 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1641
timestamp 1694700623
transform 1 0 185136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1647
timestamp 1694700623
transform 1 0 185808 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1711
timestamp 1694700623
transform 1 0 192976 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1717
timestamp 1694700623
transform 1 0 193648 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1781
timestamp 1694700623
transform 1 0 200816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1787
timestamp 1694700623
transform 1 0 201488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1803
timestamp 1694700623
transform 1 0 203280 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1811
timestamp 1694700623
transform 1 0 204176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1813
timestamp 1694700623
transform 1 0 204400 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_6
timestamp 1694700623
transform 1 0 2016 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1694700623
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1694700623
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1694700623
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1694700623
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1694700623
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1694700623
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1694700623
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1694700623
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1694700623
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1694700623
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1694700623
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1694700623
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1694700623
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1694700623
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_562
timestamp 1694700623
transform 1 0 64288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_626
timestamp 1694700623
transform 1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_632
timestamp 1694700623
transform 1 0 72128 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_696
timestamp 1694700623
transform 1 0 79296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_702
timestamp 1694700623
transform 1 0 79968 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_766
timestamp 1694700623
transform 1 0 87136 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_772
timestamp 1694700623
transform 1 0 87808 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_836
timestamp 1694700623
transform 1 0 94976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_842
timestamp 1694700623
transform 1 0 95648 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_906
timestamp 1694700623
transform 1 0 102816 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_912
timestamp 1694700623
transform 1 0 103488 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_976
timestamp 1694700623
transform 1 0 110656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_982
timestamp 1694700623
transform 1 0 111328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1046
timestamp 1694700623
transform 1 0 118496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1052
timestamp 1694700623
transform 1 0 119168 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1116
timestamp 1694700623
transform 1 0 126336 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1122
timestamp 1694700623
transform 1 0 127008 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1186
timestamp 1694700623
transform 1 0 134176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1192
timestamp 1694700623
transform 1 0 134848 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1256
timestamp 1694700623
transform 1 0 142016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1262
timestamp 1694700623
transform 1 0 142688 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1326
timestamp 1694700623
transform 1 0 149856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1332
timestamp 1694700623
transform 1 0 150528 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1396
timestamp 1694700623
transform 1 0 157696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1402
timestamp 1694700623
transform 1 0 158368 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1466
timestamp 1694700623
transform 1 0 165536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1472
timestamp 1694700623
transform 1 0 166208 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1536
timestamp 1694700623
transform 1 0 173376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1542
timestamp 1694700623
transform 1 0 174048 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1606
timestamp 1694700623
transform 1 0 181216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1612
timestamp 1694700623
transform 1 0 181888 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1676
timestamp 1694700623
transform 1 0 189056 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1682
timestamp 1694700623
transform 1 0 189728 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1746
timestamp 1694700623
transform 1 0 196896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1752
timestamp 1694700623
transform 1 0 197568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_1784
timestamp 1694700623
transform 1 0 201152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1800
timestamp 1694700623
transform 1 0 202944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1808
timestamp 1694700623
transform 1 0 203840 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1812
timestamp 1694700623
transform 1 0 204288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1694700623
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1694700623
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1694700623
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1694700623
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1694700623
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1694700623
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1694700623
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1694700623
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1694700623
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1694700623
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1694700623
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1694700623
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1694700623
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1694700623
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1694700623
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1694700623
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_527
timestamp 1694700623
transform 1 0 60368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_591
timestamp 1694700623
transform 1 0 67536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_597
timestamp 1694700623
transform 1 0 68208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_661
timestamp 1694700623
transform 1 0 75376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_667
timestamp 1694700623
transform 1 0 76048 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_731
timestamp 1694700623
transform 1 0 83216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_737
timestamp 1694700623
transform 1 0 83888 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_801
timestamp 1694700623
transform 1 0 91056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_807
timestamp 1694700623
transform 1 0 91728 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_871
timestamp 1694700623
transform 1 0 98896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_877
timestamp 1694700623
transform 1 0 99568 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_941
timestamp 1694700623
transform 1 0 106736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_947
timestamp 1694700623
transform 1 0 107408 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1011
timestamp 1694700623
transform 1 0 114576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1017
timestamp 1694700623
transform 1 0 115248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1081
timestamp 1694700623
transform 1 0 122416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1087
timestamp 1694700623
transform 1 0 123088 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1151
timestamp 1694700623
transform 1 0 130256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1157
timestamp 1694700623
transform 1 0 130928 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1221
timestamp 1694700623
transform 1 0 138096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1227
timestamp 1694700623
transform 1 0 138768 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1291
timestamp 1694700623
transform 1 0 145936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1297
timestamp 1694700623
transform 1 0 146608 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1361
timestamp 1694700623
transform 1 0 153776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1367
timestamp 1694700623
transform 1 0 154448 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1431
timestamp 1694700623
transform 1 0 161616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1437
timestamp 1694700623
transform 1 0 162288 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1501
timestamp 1694700623
transform 1 0 169456 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1507
timestamp 1694700623
transform 1 0 170128 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1571
timestamp 1694700623
transform 1 0 177296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1577
timestamp 1694700623
transform 1 0 177968 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1641
timestamp 1694700623
transform 1 0 185136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1647
timestamp 1694700623
transform 1 0 185808 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1711
timestamp 1694700623
transform 1 0 192976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1717
timestamp 1694700623
transform 1 0 193648 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1781
timestamp 1694700623
transform 1 0 200816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1787
timestamp 1694700623
transform 1 0 201488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1803
timestamp 1694700623
transform 1 0 203280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1811
timestamp 1694700623
transform 1 0 204176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1813
timestamp 1694700623
transform 1 0 204400 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1694700623
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1694700623
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1694700623
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1694700623
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1694700623
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1694700623
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1694700623
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1694700623
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1694700623
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1694700623
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1694700623
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1694700623
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1694700623
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1694700623
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1694700623
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1694700623
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_562
timestamp 1694700623
transform 1 0 64288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_626
timestamp 1694700623
transform 1 0 71456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_632
timestamp 1694700623
transform 1 0 72128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_696
timestamp 1694700623
transform 1 0 79296 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_702
timestamp 1694700623
transform 1 0 79968 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_766
timestamp 1694700623
transform 1 0 87136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_772
timestamp 1694700623
transform 1 0 87808 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_836
timestamp 1694700623
transform 1 0 94976 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_842
timestamp 1694700623
transform 1 0 95648 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_906
timestamp 1694700623
transform 1 0 102816 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_912
timestamp 1694700623
transform 1 0 103488 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_976
timestamp 1694700623
transform 1 0 110656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_982
timestamp 1694700623
transform 1 0 111328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1046
timestamp 1694700623
transform 1 0 118496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1052
timestamp 1694700623
transform 1 0 119168 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1116
timestamp 1694700623
transform 1 0 126336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1122
timestamp 1694700623
transform 1 0 127008 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1186
timestamp 1694700623
transform 1 0 134176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1192
timestamp 1694700623
transform 1 0 134848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1256
timestamp 1694700623
transform 1 0 142016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1262
timestamp 1694700623
transform 1 0 142688 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1326
timestamp 1694700623
transform 1 0 149856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1332
timestamp 1694700623
transform 1 0 150528 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1396
timestamp 1694700623
transform 1 0 157696 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1402
timestamp 1694700623
transform 1 0 158368 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1466
timestamp 1694700623
transform 1 0 165536 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1472
timestamp 1694700623
transform 1 0 166208 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1536
timestamp 1694700623
transform 1 0 173376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1542
timestamp 1694700623
transform 1 0 174048 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1606
timestamp 1694700623
transform 1 0 181216 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1612
timestamp 1694700623
transform 1 0 181888 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1676
timestamp 1694700623
transform 1 0 189056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1682
timestamp 1694700623
transform 1 0 189728 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1746
timestamp 1694700623
transform 1 0 196896 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_1752
timestamp 1694700623
transform 1 0 197568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1784
timestamp 1694700623
transform 1 0 201152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1800
timestamp 1694700623
transform 1 0 202944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1808
timestamp 1694700623
transform 1 0 203840 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1812
timestamp 1694700623
transform 1 0 204288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1694700623
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1694700623
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1694700623
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1694700623
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1694700623
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1694700623
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1694700623
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1694700623
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1694700623
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1694700623
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1694700623
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1694700623
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1694700623
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1694700623
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1694700623
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1694700623
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1694700623
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1694700623
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_597
timestamp 1694700623
transform 1 0 68208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_661
timestamp 1694700623
transform 1 0 75376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_667
timestamp 1694700623
transform 1 0 76048 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_731
timestamp 1694700623
transform 1 0 83216 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_737
timestamp 1694700623
transform 1 0 83888 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_801
timestamp 1694700623
transform 1 0 91056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_807
timestamp 1694700623
transform 1 0 91728 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_871
timestamp 1694700623
transform 1 0 98896 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_877
timestamp 1694700623
transform 1 0 99568 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_941
timestamp 1694700623
transform 1 0 106736 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_947
timestamp 1694700623
transform 1 0 107408 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1011
timestamp 1694700623
transform 1 0 114576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1017
timestamp 1694700623
transform 1 0 115248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1081
timestamp 1694700623
transform 1 0 122416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1087
timestamp 1694700623
transform 1 0 123088 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1151
timestamp 1694700623
transform 1 0 130256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1157
timestamp 1694700623
transform 1 0 130928 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1221
timestamp 1694700623
transform 1 0 138096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1227
timestamp 1694700623
transform 1 0 138768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1291
timestamp 1694700623
transform 1 0 145936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1297
timestamp 1694700623
transform 1 0 146608 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1361
timestamp 1694700623
transform 1 0 153776 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1367
timestamp 1694700623
transform 1 0 154448 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1431
timestamp 1694700623
transform 1 0 161616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1437
timestamp 1694700623
transform 1 0 162288 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1501
timestamp 1694700623
transform 1 0 169456 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1507
timestamp 1694700623
transform 1 0 170128 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1571
timestamp 1694700623
transform 1 0 177296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1577
timestamp 1694700623
transform 1 0 177968 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1641
timestamp 1694700623
transform 1 0 185136 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1647
timestamp 1694700623
transform 1 0 185808 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1711
timestamp 1694700623
transform 1 0 192976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1717
timestamp 1694700623
transform 1 0 193648 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1781
timestamp 1694700623
transform 1 0 200816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1787
timestamp 1694700623
transform 1 0 201488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1803
timestamp 1694700623
transform 1 0 203280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1811
timestamp 1694700623
transform 1 0 204176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1813
timestamp 1694700623
transform 1 0 204400 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1694700623
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1694700623
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1694700623
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1694700623
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1694700623
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1694700623
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1694700623
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1694700623
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1694700623
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1694700623
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1694700623
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1694700623
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1694700623
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1694700623
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1694700623
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1694700623
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1694700623
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1694700623
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_632
timestamp 1694700623
transform 1 0 72128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_696
timestamp 1694700623
transform 1 0 79296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_702
timestamp 1694700623
transform 1 0 79968 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_766
timestamp 1694700623
transform 1 0 87136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_772
timestamp 1694700623
transform 1 0 87808 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_836
timestamp 1694700623
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_842
timestamp 1694700623
transform 1 0 95648 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_906
timestamp 1694700623
transform 1 0 102816 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_912
timestamp 1694700623
transform 1 0 103488 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_976
timestamp 1694700623
transform 1 0 110656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_982
timestamp 1694700623
transform 1 0 111328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1046
timestamp 1694700623
transform 1 0 118496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1052
timestamp 1694700623
transform 1 0 119168 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1116
timestamp 1694700623
transform 1 0 126336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1122
timestamp 1694700623
transform 1 0 127008 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1186
timestamp 1694700623
transform 1 0 134176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1192
timestamp 1694700623
transform 1 0 134848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1256
timestamp 1694700623
transform 1 0 142016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1262
timestamp 1694700623
transform 1 0 142688 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1326
timestamp 1694700623
transform 1 0 149856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1332
timestamp 1694700623
transform 1 0 150528 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1396
timestamp 1694700623
transform 1 0 157696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1402
timestamp 1694700623
transform 1 0 158368 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1466
timestamp 1694700623
transform 1 0 165536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1472
timestamp 1694700623
transform 1 0 166208 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1536
timestamp 1694700623
transform 1 0 173376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1542
timestamp 1694700623
transform 1 0 174048 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1606
timestamp 1694700623
transform 1 0 181216 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1612
timestamp 1694700623
transform 1 0 181888 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1676
timestamp 1694700623
transform 1 0 189056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1682
timestamp 1694700623
transform 1 0 189728 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1746
timestamp 1694700623
transform 1 0 196896 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_1752
timestamp 1694700623
transform 1 0 197568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1784
timestamp 1694700623
transform 1 0 201152 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1800
timestamp 1694700623
transform 1 0 202944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1808
timestamp 1694700623
transform 1 0 203840 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1812
timestamp 1694700623
transform 1 0 204288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1694700623
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1694700623
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1694700623
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1694700623
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1694700623
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1694700623
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1694700623
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1694700623
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1694700623
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1694700623
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1694700623
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1694700623
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1694700623
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1694700623
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1694700623
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1694700623
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1694700623
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1694700623
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1694700623
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1694700623
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1694700623
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_597
timestamp 1694700623
transform 1 0 68208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_661
timestamp 1694700623
transform 1 0 75376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_667
timestamp 1694700623
transform 1 0 76048 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_731
timestamp 1694700623
transform 1 0 83216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_737
timestamp 1694700623
transform 1 0 83888 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_801
timestamp 1694700623
transform 1 0 91056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_807
timestamp 1694700623
transform 1 0 91728 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_871
timestamp 1694700623
transform 1 0 98896 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_877
timestamp 1694700623
transform 1 0 99568 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_941
timestamp 1694700623
transform 1 0 106736 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_947
timestamp 1694700623
transform 1 0 107408 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1011
timestamp 1694700623
transform 1 0 114576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1017
timestamp 1694700623
transform 1 0 115248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1081
timestamp 1694700623
transform 1 0 122416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1087
timestamp 1694700623
transform 1 0 123088 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1151
timestamp 1694700623
transform 1 0 130256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1157
timestamp 1694700623
transform 1 0 130928 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1221
timestamp 1694700623
transform 1 0 138096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1227
timestamp 1694700623
transform 1 0 138768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1291
timestamp 1694700623
transform 1 0 145936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1297
timestamp 1694700623
transform 1 0 146608 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1361
timestamp 1694700623
transform 1 0 153776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1367
timestamp 1694700623
transform 1 0 154448 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1431
timestamp 1694700623
transform 1 0 161616 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1437
timestamp 1694700623
transform 1 0 162288 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1501
timestamp 1694700623
transform 1 0 169456 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1507
timestamp 1694700623
transform 1 0 170128 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1571
timestamp 1694700623
transform 1 0 177296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1577
timestamp 1694700623
transform 1 0 177968 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1641
timestamp 1694700623
transform 1 0 185136 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1647
timestamp 1694700623
transform 1 0 185808 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1711
timestamp 1694700623
transform 1 0 192976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1717
timestamp 1694700623
transform 1 0 193648 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1781
timestamp 1694700623
transform 1 0 200816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_1787
timestamp 1694700623
transform 1 0 201488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1803
timestamp 1694700623
transform 1 0 203280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1811
timestamp 1694700623
transform 1 0 204176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1813
timestamp 1694700623
transform 1 0 204400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1694700623
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1694700623
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1694700623
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1694700623
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1694700623
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1694700623
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1694700623
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1694700623
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1694700623
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1694700623
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1694700623
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1694700623
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1694700623
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1694700623
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1694700623
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1694700623
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1694700623
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1694700623
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_632
timestamp 1694700623
transform 1 0 72128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_696
timestamp 1694700623
transform 1 0 79296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_702
timestamp 1694700623
transform 1 0 79968 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_766
timestamp 1694700623
transform 1 0 87136 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_772
timestamp 1694700623
transform 1 0 87808 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_836
timestamp 1694700623
transform 1 0 94976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_842
timestamp 1694700623
transform 1 0 95648 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_906
timestamp 1694700623
transform 1 0 102816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_912
timestamp 1694700623
transform 1 0 103488 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_976
timestamp 1694700623
transform 1 0 110656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_982
timestamp 1694700623
transform 1 0 111328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1046
timestamp 1694700623
transform 1 0 118496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1052
timestamp 1694700623
transform 1 0 119168 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1116
timestamp 1694700623
transform 1 0 126336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1122
timestamp 1694700623
transform 1 0 127008 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1186
timestamp 1694700623
transform 1 0 134176 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1192
timestamp 1694700623
transform 1 0 134848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1256
timestamp 1694700623
transform 1 0 142016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1262
timestamp 1694700623
transform 1 0 142688 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1326
timestamp 1694700623
transform 1 0 149856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1332
timestamp 1694700623
transform 1 0 150528 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1396
timestamp 1694700623
transform 1 0 157696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1402
timestamp 1694700623
transform 1 0 158368 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1466
timestamp 1694700623
transform 1 0 165536 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1472
timestamp 1694700623
transform 1 0 166208 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1536
timestamp 1694700623
transform 1 0 173376 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1542
timestamp 1694700623
transform 1 0 174048 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1606
timestamp 1694700623
transform 1 0 181216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1612
timestamp 1694700623
transform 1 0 181888 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1676
timestamp 1694700623
transform 1 0 189056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1682
timestamp 1694700623
transform 1 0 189728 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1746
timestamp 1694700623
transform 1 0 196896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_1752
timestamp 1694700623
transform 1 0 197568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_1784
timestamp 1694700623
transform 1 0 201152 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1800
timestamp 1694700623
transform 1 0 202944 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1808
timestamp 1694700623
transform 1 0 203840 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1812
timestamp 1694700623
transform 1 0 204288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1694700623
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1694700623
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1694700623
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1694700623
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1694700623
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1694700623
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1694700623
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1694700623
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1694700623
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1694700623
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1694700623
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1694700623
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1694700623
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1694700623
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1694700623
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1694700623
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1694700623
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1694700623
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1694700623
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1694700623
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_667
timestamp 1694700623
transform 1 0 76048 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_731
timestamp 1694700623
transform 1 0 83216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_737
timestamp 1694700623
transform 1 0 83888 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_801
timestamp 1694700623
transform 1 0 91056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_807
timestamp 1694700623
transform 1 0 91728 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_871
timestamp 1694700623
transform 1 0 98896 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_877
timestamp 1694700623
transform 1 0 99568 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_941
timestamp 1694700623
transform 1 0 106736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_947
timestamp 1694700623
transform 1 0 107408 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1011
timestamp 1694700623
transform 1 0 114576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1017
timestamp 1694700623
transform 1 0 115248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1081
timestamp 1694700623
transform 1 0 122416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1087
timestamp 1694700623
transform 1 0 123088 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1151
timestamp 1694700623
transform 1 0 130256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1157
timestamp 1694700623
transform 1 0 130928 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1221
timestamp 1694700623
transform 1 0 138096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1227
timestamp 1694700623
transform 1 0 138768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1291
timestamp 1694700623
transform 1 0 145936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1297
timestamp 1694700623
transform 1 0 146608 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1361
timestamp 1694700623
transform 1 0 153776 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1367
timestamp 1694700623
transform 1 0 154448 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1431
timestamp 1694700623
transform 1 0 161616 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1437
timestamp 1694700623
transform 1 0 162288 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1501
timestamp 1694700623
transform 1 0 169456 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1507
timestamp 1694700623
transform 1 0 170128 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1571
timestamp 1694700623
transform 1 0 177296 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1577
timestamp 1694700623
transform 1 0 177968 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1641
timestamp 1694700623
transform 1 0 185136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1647
timestamp 1694700623
transform 1 0 185808 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1711
timestamp 1694700623
transform 1 0 192976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1717
timestamp 1694700623
transform 1 0 193648 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1781
timestamp 1694700623
transform 1 0 200816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_1787
timestamp 1694700623
transform 1 0 201488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_1803
timestamp 1694700623
transform 1 0 203280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1811
timestamp 1694700623
transform 1 0 204176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1813
timestamp 1694700623
transform 1 0 204400 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1694700623
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1694700623
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1694700623
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1694700623
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1694700623
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1694700623
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1694700623
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1694700623
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1694700623
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1694700623
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1694700623
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1694700623
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1694700623
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1694700623
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1694700623
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1694700623
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1694700623
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1694700623
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_632
timestamp 1694700623
transform 1 0 72128 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_696
timestamp 1694700623
transform 1 0 79296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_702
timestamp 1694700623
transform 1 0 79968 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_766
timestamp 1694700623
transform 1 0 87136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_772
timestamp 1694700623
transform 1 0 87808 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_836
timestamp 1694700623
transform 1 0 94976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_842
timestamp 1694700623
transform 1 0 95648 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_906
timestamp 1694700623
transform 1 0 102816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_912
timestamp 1694700623
transform 1 0 103488 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_976
timestamp 1694700623
transform 1 0 110656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_982
timestamp 1694700623
transform 1 0 111328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1046
timestamp 1694700623
transform 1 0 118496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1052
timestamp 1694700623
transform 1 0 119168 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1116
timestamp 1694700623
transform 1 0 126336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1122
timestamp 1694700623
transform 1 0 127008 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1186
timestamp 1694700623
transform 1 0 134176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1192
timestamp 1694700623
transform 1 0 134848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1256
timestamp 1694700623
transform 1 0 142016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1262
timestamp 1694700623
transform 1 0 142688 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1326
timestamp 1694700623
transform 1 0 149856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1332
timestamp 1694700623
transform 1 0 150528 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1396
timestamp 1694700623
transform 1 0 157696 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1402
timestamp 1694700623
transform 1 0 158368 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1466
timestamp 1694700623
transform 1 0 165536 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1472
timestamp 1694700623
transform 1 0 166208 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1536
timestamp 1694700623
transform 1 0 173376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1542
timestamp 1694700623
transform 1 0 174048 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1606
timestamp 1694700623
transform 1 0 181216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1612
timestamp 1694700623
transform 1 0 181888 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1676
timestamp 1694700623
transform 1 0 189056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1682
timestamp 1694700623
transform 1 0 189728 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1746
timestamp 1694700623
transform 1 0 196896 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_1752
timestamp 1694700623
transform 1 0 197568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_1784
timestamp 1694700623
transform 1 0 201152 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1800
timestamp 1694700623
transform 1 0 202944 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1808
timestamp 1694700623
transform 1 0 203840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_1812
timestamp 1694700623
transform 1 0 204288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1694700623
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1694700623
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1694700623
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1694700623
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1694700623
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1694700623
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1694700623
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1694700623
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1694700623
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1694700623
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1694700623
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1694700623
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1694700623
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1694700623
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1694700623
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1694700623
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1694700623
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1694700623
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1694700623
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1694700623
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_667
timestamp 1694700623
transform 1 0 76048 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_731
timestamp 1694700623
transform 1 0 83216 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_737
timestamp 1694700623
transform 1 0 83888 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_801
timestamp 1694700623
transform 1 0 91056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_807
timestamp 1694700623
transform 1 0 91728 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_871
timestamp 1694700623
transform 1 0 98896 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_877
timestamp 1694700623
transform 1 0 99568 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_941
timestamp 1694700623
transform 1 0 106736 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_947
timestamp 1694700623
transform 1 0 107408 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1011
timestamp 1694700623
transform 1 0 114576 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1017
timestamp 1694700623
transform 1 0 115248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1081
timestamp 1694700623
transform 1 0 122416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1087
timestamp 1694700623
transform 1 0 123088 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1151
timestamp 1694700623
transform 1 0 130256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1157
timestamp 1694700623
transform 1 0 130928 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1221
timestamp 1694700623
transform 1 0 138096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1227
timestamp 1694700623
transform 1 0 138768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1291
timestamp 1694700623
transform 1 0 145936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1297
timestamp 1694700623
transform 1 0 146608 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1361
timestamp 1694700623
transform 1 0 153776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1367
timestamp 1694700623
transform 1 0 154448 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1431
timestamp 1694700623
transform 1 0 161616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1437
timestamp 1694700623
transform 1 0 162288 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1501
timestamp 1694700623
transform 1 0 169456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1507
timestamp 1694700623
transform 1 0 170128 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1571
timestamp 1694700623
transform 1 0 177296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1577
timestamp 1694700623
transform 1 0 177968 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1641
timestamp 1694700623
transform 1 0 185136 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1647
timestamp 1694700623
transform 1 0 185808 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1711
timestamp 1694700623
transform 1 0 192976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1717
timestamp 1694700623
transform 1 0 193648 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1781
timestamp 1694700623
transform 1 0 200816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_1787
timestamp 1694700623
transform 1 0 201488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_1803
timestamp 1694700623
transform 1 0 203280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_1811
timestamp 1694700623
transform 1 0 204176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_1813
timestamp 1694700623
transform 1 0 204400 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_6
timestamp 1694700623
transform 1 0 2016 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1694700623
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1694700623
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1694700623
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1694700623
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1694700623
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1694700623
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1694700623
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1694700623
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1694700623
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1694700623
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1694700623
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1694700623
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1694700623
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1694700623
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1694700623
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1694700623
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_632
timestamp 1694700623
transform 1 0 72128 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_696
timestamp 1694700623
transform 1 0 79296 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_702
timestamp 1694700623
transform 1 0 79968 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_766
timestamp 1694700623
transform 1 0 87136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_772
timestamp 1694700623
transform 1 0 87808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_836
timestamp 1694700623
transform 1 0 94976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_842
timestamp 1694700623
transform 1 0 95648 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_906
timestamp 1694700623
transform 1 0 102816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_912
timestamp 1694700623
transform 1 0 103488 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_976
timestamp 1694700623
transform 1 0 110656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_982
timestamp 1694700623
transform 1 0 111328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1046
timestamp 1694700623
transform 1 0 118496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1052
timestamp 1694700623
transform 1 0 119168 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1116
timestamp 1694700623
transform 1 0 126336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1122
timestamp 1694700623
transform 1 0 127008 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1186
timestamp 1694700623
transform 1 0 134176 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1192
timestamp 1694700623
transform 1 0 134848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1256
timestamp 1694700623
transform 1 0 142016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1262
timestamp 1694700623
transform 1 0 142688 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1326
timestamp 1694700623
transform 1 0 149856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1332
timestamp 1694700623
transform 1 0 150528 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1396
timestamp 1694700623
transform 1 0 157696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1402
timestamp 1694700623
transform 1 0 158368 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1466
timestamp 1694700623
transform 1 0 165536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1472
timestamp 1694700623
transform 1 0 166208 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1536
timestamp 1694700623
transform 1 0 173376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1542
timestamp 1694700623
transform 1 0 174048 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1606
timestamp 1694700623
transform 1 0 181216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1612
timestamp 1694700623
transform 1 0 181888 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1676
timestamp 1694700623
transform 1 0 189056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1682
timestamp 1694700623
transform 1 0 189728 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1746
timestamp 1694700623
transform 1 0 196896 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_1752
timestamp 1694700623
transform 1 0 197568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_1784
timestamp 1694700623
transform 1 0 201152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_1800
timestamp 1694700623
transform 1 0 202944 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1808
timestamp 1694700623
transform 1 0 203840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1694700623
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1694700623
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1694700623
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1694700623
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1694700623
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1694700623
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1694700623
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1694700623
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1694700623
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1694700623
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1694700623
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1694700623
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1694700623
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1694700623
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1694700623
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1694700623
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1694700623
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1694700623
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1694700623
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1694700623
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_667
timestamp 1694700623
transform 1 0 76048 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_731
timestamp 1694700623
transform 1 0 83216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_737
timestamp 1694700623
transform 1 0 83888 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_801
timestamp 1694700623
transform 1 0 91056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_807
timestamp 1694700623
transform 1 0 91728 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_871
timestamp 1694700623
transform 1 0 98896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_877
timestamp 1694700623
transform 1 0 99568 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_941
timestamp 1694700623
transform 1 0 106736 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_947
timestamp 1694700623
transform 1 0 107408 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1011
timestamp 1694700623
transform 1 0 114576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1017
timestamp 1694700623
transform 1 0 115248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1081
timestamp 1694700623
transform 1 0 122416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1087
timestamp 1694700623
transform 1 0 123088 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1151
timestamp 1694700623
transform 1 0 130256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1157
timestamp 1694700623
transform 1 0 130928 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1221
timestamp 1694700623
transform 1 0 138096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1227
timestamp 1694700623
transform 1 0 138768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1291
timestamp 1694700623
transform 1 0 145936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1297
timestamp 1694700623
transform 1 0 146608 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1361
timestamp 1694700623
transform 1 0 153776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1367
timestamp 1694700623
transform 1 0 154448 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1431
timestamp 1694700623
transform 1 0 161616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1437
timestamp 1694700623
transform 1 0 162288 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1501
timestamp 1694700623
transform 1 0 169456 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1507
timestamp 1694700623
transform 1 0 170128 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1571
timestamp 1694700623
transform 1 0 177296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1577
timestamp 1694700623
transform 1 0 177968 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1641
timestamp 1694700623
transform 1 0 185136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1647
timestamp 1694700623
transform 1 0 185808 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1711
timestamp 1694700623
transform 1 0 192976 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1717
timestamp 1694700623
transform 1 0 193648 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1781
timestamp 1694700623
transform 1 0 200816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_1787
timestamp 1694700623
transform 1 0 201488 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1694700623
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1694700623
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1694700623
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1694700623
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1694700623
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1694700623
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1694700623
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1694700623
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1694700623
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1694700623
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1694700623
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1694700623
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1694700623
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1694700623
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1694700623
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1694700623
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1694700623
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1694700623
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_632
timestamp 1694700623
transform 1 0 72128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_696
timestamp 1694700623
transform 1 0 79296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_702
timestamp 1694700623
transform 1 0 79968 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_766
timestamp 1694700623
transform 1 0 87136 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_772
timestamp 1694700623
transform 1 0 87808 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_836
timestamp 1694700623
transform 1 0 94976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_842
timestamp 1694700623
transform 1 0 95648 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_906
timestamp 1694700623
transform 1 0 102816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_912
timestamp 1694700623
transform 1 0 103488 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_976
timestamp 1694700623
transform 1 0 110656 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_982
timestamp 1694700623
transform 1 0 111328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1046
timestamp 1694700623
transform 1 0 118496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1052
timestamp 1694700623
transform 1 0 119168 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1116
timestamp 1694700623
transform 1 0 126336 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1122
timestamp 1694700623
transform 1 0 127008 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1186
timestamp 1694700623
transform 1 0 134176 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1192
timestamp 1694700623
transform 1 0 134848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1256
timestamp 1694700623
transform 1 0 142016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1262
timestamp 1694700623
transform 1 0 142688 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1326
timestamp 1694700623
transform 1 0 149856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1332
timestamp 1694700623
transform 1 0 150528 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1396
timestamp 1694700623
transform 1 0 157696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1402
timestamp 1694700623
transform 1 0 158368 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1466
timestamp 1694700623
transform 1 0 165536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1472
timestamp 1694700623
transform 1 0 166208 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1536
timestamp 1694700623
transform 1 0 173376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1542
timestamp 1694700623
transform 1 0 174048 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1606
timestamp 1694700623
transform 1 0 181216 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1612
timestamp 1694700623
transform 1 0 181888 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1676
timestamp 1694700623
transform 1 0 189056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1682
timestamp 1694700623
transform 1 0 189728 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1746
timestamp 1694700623
transform 1 0 196896 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_1752
timestamp 1694700623
transform 1 0 197568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_1784
timestamp 1694700623
transform 1 0 201152 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_1800
timestamp 1694700623
transform 1 0 202944 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1808
timestamp 1694700623
transform 1 0 203840 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_1812
timestamp 1694700623
transform 1 0 204288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1694700623
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1694700623
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1694700623
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1694700623
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1694700623
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1694700623
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1694700623
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1694700623
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1694700623
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1694700623
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1694700623
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1694700623
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1694700623
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1694700623
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1694700623
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1694700623
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1694700623
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1694700623
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1694700623
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1694700623
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_667
timestamp 1694700623
transform 1 0 76048 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_731
timestamp 1694700623
transform 1 0 83216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_737
timestamp 1694700623
transform 1 0 83888 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_801
timestamp 1694700623
transform 1 0 91056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_807
timestamp 1694700623
transform 1 0 91728 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_871
timestamp 1694700623
transform 1 0 98896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_877
timestamp 1694700623
transform 1 0 99568 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_941
timestamp 1694700623
transform 1 0 106736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_947
timestamp 1694700623
transform 1 0 107408 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1011
timestamp 1694700623
transform 1 0 114576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1017
timestamp 1694700623
transform 1 0 115248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1081
timestamp 1694700623
transform 1 0 122416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1087
timestamp 1694700623
transform 1 0 123088 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1151
timestamp 1694700623
transform 1 0 130256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1157
timestamp 1694700623
transform 1 0 130928 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1221
timestamp 1694700623
transform 1 0 138096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1227
timestamp 1694700623
transform 1 0 138768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1291
timestamp 1694700623
transform 1 0 145936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1297
timestamp 1694700623
transform 1 0 146608 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1361
timestamp 1694700623
transform 1 0 153776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1367
timestamp 1694700623
transform 1 0 154448 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1431
timestamp 1694700623
transform 1 0 161616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1437
timestamp 1694700623
transform 1 0 162288 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1501
timestamp 1694700623
transform 1 0 169456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1507
timestamp 1694700623
transform 1 0 170128 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1571
timestamp 1694700623
transform 1 0 177296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1577
timestamp 1694700623
transform 1 0 177968 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1641
timestamp 1694700623
transform 1 0 185136 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1647
timestamp 1694700623
transform 1 0 185808 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1711
timestamp 1694700623
transform 1 0 192976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1717
timestamp 1694700623
transform 1 0 193648 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1781
timestamp 1694700623
transform 1 0 200816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_1787
timestamp 1694700623
transform 1 0 201488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_1803
timestamp 1694700623
transform 1 0 203280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_1811
timestamp 1694700623
transform 1 0 204176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_1813
timestamp 1694700623
transform 1 0 204400 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1694700623
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_36
timestamp 1694700623
transform 1 0 5376 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_70
timestamp 1694700623
transform 1 0 9184 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_104
timestamp 1694700623
transform 1 0 12992 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_138
timestamp 1694700623
transform 1 0 16800 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_172
timestamp 1694700623
transform 1 0 20608 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_206
timestamp 1694700623
transform 1 0 24416 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_240
timestamp 1694700623
transform 1 0 28224 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_274
timestamp 1694700623
transform 1 0 32032 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_308
timestamp 1694700623
transform 1 0 35840 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_342
timestamp 1694700623
transform 1 0 39648 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_376
timestamp 1694700623
transform 1 0 43456 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_384
timestamp 1694700623
transform 1 0 44352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_386
timestamp 1694700623
transform 1 0 44576 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_389
timestamp 1694700623
transform 1 0 44912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_405
timestamp 1694700623
transform 1 0 46704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_407
timestamp 1694700623
transform 1 0 46928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_410
timestamp 1694700623
transform 1 0 47264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_420
timestamp 1694700623
transform 1 0 48384 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_436
timestamp 1694700623
transform 1 0 50176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_440
timestamp 1694700623
transform 1 0 50624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_444
timestamp 1694700623
transform 1 0 51072 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_450
timestamp 1694700623
transform 1 0 51744 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_466
timestamp 1694700623
transform 1 0 53536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_474
timestamp 1694700623
transform 1 0 54432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_478
timestamp 1694700623
transform 1 0 54880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_482
timestamp 1694700623
transform 1 0 55328 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_498
timestamp 1694700623
transform 1 0 57120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_506
timestamp 1694700623
transform 1 0 58016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_512
timestamp 1694700623
transform 1 0 58688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_516
timestamp 1694700623
transform 1 0 59136 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_532
timestamp 1694700623
transform 1 0 60928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_542
timestamp 1694700623
transform 1 0 62048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_546
timestamp 1694700623
transform 1 0 62496 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_562
timestamp 1694700623
transform 1 0 64288 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_570
timestamp 1694700623
transform 1 0 65184 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_573
timestamp 1694700623
transform 1 0 65520 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_577
timestamp 1694700623
transform 1 0 65968 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_580
timestamp 1694700623
transform 1 0 66304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_588
timestamp 1694700623
transform 1 0 67200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_592
timestamp 1694700623
transform 1 0 67648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_596
timestamp 1694700623
transform 1 0 68096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_600
timestamp 1694700623
transform 1 0 68544 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_603
timestamp 1694700623
transform 1 0 68880 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_611
timestamp 1694700623
transform 1 0 69776 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_614
timestamp 1694700623
transform 1 0 70112 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_630
timestamp 1694700623
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_634
timestamp 1694700623
transform 1 0 72352 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_642
timestamp 1694700623
transform 1 0 73248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_648
timestamp 1694700623
transform 1 0 73920 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_656
timestamp 1694700623
transform 1 0 74816 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_660
timestamp 1694700623
transform 1 0 75264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_664
timestamp 1694700623
transform 1 0 75712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_682
timestamp 1694700623
transform 1 0 77728 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_690
timestamp 1694700623
transform 1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_692
timestamp 1694700623
transform 1 0 78848 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_695
timestamp 1694700623
transform 1 0 79184 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_711
timestamp 1694700623
transform 1 0 80976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_713
timestamp 1694700623
transform 1 0 81200 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_716
timestamp 1694700623
transform 1 0 81536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_720
timestamp 1694700623
transform 1 0 81984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_722
timestamp 1694700623
transform 1 0 82208 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_725
timestamp 1694700623
transform 1 0 82544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_729
timestamp 1694700623
transform 1 0 82992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_745
timestamp 1694700623
transform 1 0 84784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_747
timestamp 1694700623
transform 1 0 85008 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_750
timestamp 1694700623
transform 1 0 85344 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_784
timestamp 1694700623
transform 1 0 89152 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_818
timestamp 1694700623
transform 1 0 92960 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_852
timestamp 1694700623
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_856
timestamp 1694700623
transform 1 0 97216 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_872
timestamp 1694700623
transform 1 0 99008 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_880
timestamp 1694700623
transform 1 0 99904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_886
timestamp 1694700623
transform 1 0 100576 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_920
timestamp 1694700623
transform 1 0 104384 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_954
timestamp 1694700623
transform 1 0 108192 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_970
timestamp 1694700623
transform 1 0 109984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_978
timestamp 1694700623
transform 1 0 110880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_982
timestamp 1694700623
transform 1 0 111328 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_988
timestamp 1694700623
transform 1 0 112000 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1022
timestamp 1694700623
transform 1 0 115808 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1056
timestamp 1694700623
transform 1 0 119616 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_1090
timestamp 1694700623
transform 1 0 123424 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1106
timestamp 1694700623
transform 1 0 125216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1110
timestamp 1694700623
transform 1 0 125664 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1118
timestamp 1694700623
transform 1 0 126560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1124
timestamp 1694700623
transform 1 0 127232 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1158
timestamp 1694700623
transform 1 0 131040 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1192
timestamp 1694700623
transform 1 0 134848 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1226
timestamp 1694700623
transform 1 0 138656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1234
timestamp 1694700623
transform 1 0 139552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_1236
timestamp 1694700623
transform 1 0 139776 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_1239
timestamp 1694700623
transform 1 0 140112 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1255
timestamp 1694700623
transform 1 0 141904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_1257
timestamp 1694700623
transform 1 0 142128 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1260
timestamp 1694700623
transform 1 0 142464 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1294
timestamp 1694700623
transform 1 0 146272 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1328
timestamp 1694700623
transform 1 0 150080 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1362
timestamp 1694700623
transform 1 0 153888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_1364
timestamp 1694700623
transform 1 0 154112 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_1367
timestamp 1694700623
transform 1 0 154448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1383
timestamp 1694700623
transform 1 0 156240 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1391
timestamp 1694700623
transform 1 0 157136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_1393
timestamp 1694700623
transform 1 0 157360 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1396
timestamp 1694700623
transform 1 0 157696 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1430
timestamp 1694700623
transform 1 0 161504 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1464
timestamp 1694700623
transform 1 0 165312 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1498
timestamp 1694700623
transform 1 0 169120 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1532
timestamp 1694700623
transform 1 0 172928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1566
timestamp 1694700623
transform 1 0 176736 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1600
timestamp 1694700623
transform 1 0 180544 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1634
timestamp 1694700623
transform 1 0 184352 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1668
timestamp 1694700623
transform 1 0 188160 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1702
timestamp 1694700623
transform 1 0 191968 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1736
timestamp 1694700623
transform 1 0 195776 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1770
timestamp 1694700623
transform 1 0 199584 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1804
timestamp 1694700623
transform 1 0 203392 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1812
timestamp 1694700623
transform 1 0 204288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_6
timestamp 1694700623
transform 1 0 2016 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_22
timestamp 1694700623
transform 1 0 3808 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_30
timestamp 1694700623
transform 1 0 4704 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1694700623
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1694700623
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1694700623
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1694700623
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_139
timestamp 1694700623
transform 1 0 16912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_143
timestamp 1694700623
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_145
timestamp 1694700623
transform 1 0 17584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_1671
timestamp 1694700623
transform 1 0 188496 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_1703
timestamp 1694700623
transform 1 0 192080 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1706
timestamp 1694700623
transform 1 0 192416 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1770
timestamp 1694700623
transform 1 0 199584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_1776
timestamp 1694700623
transform 1 0 200256 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1808
timestamp 1694700623
transform 1 0 203840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_1812
timestamp 1694700623
transform 1 0 204288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1694700623
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1694700623
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1694700623
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1694700623
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1694700623
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1671
timestamp 1694700623
transform 1 0 188496 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1735
timestamp 1694700623
transform 1 0 195664 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1741
timestamp 1694700623
transform 1 0 196336 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1805
timestamp 1694700623
transform 1 0 203504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_1811
timestamp 1694700623
transform 1 0 204176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_1813
timestamp 1694700623
transform 1 0 204400 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1694700623
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1694700623
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1694700623
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1694700623
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_107
timestamp 1694700623
transform 1 0 13328 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_139
timestamp 1694700623
transform 1 0 16912 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_143
timestamp 1694700623
transform 1 0 17360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_145
timestamp 1694700623
transform 1 0 17584 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_1671
timestamp 1694700623
transform 1 0 188496 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_1703
timestamp 1694700623
transform 1 0 192080 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1706
timestamp 1694700623
transform 1 0 192416 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1770
timestamp 1694700623
transform 1 0 199584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_1776
timestamp 1694700623
transform 1 0 200256 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1808
timestamp 1694700623
transform 1 0 203840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_1812
timestamp 1694700623
transform 1 0 204288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1694700623
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1694700623
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1694700623
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1694700623
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1694700623
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1671
timestamp 1694700623
transform 1 0 188496 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1735
timestamp 1694700623
transform 1 0 195664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1741
timestamp 1694700623
transform 1 0 196336 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1805
timestamp 1694700623
transform 1 0 203504 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_1811
timestamp 1694700623
transform 1 0 204176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_1813
timestamp 1694700623
transform 1 0 204400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1694700623
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1694700623
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1694700623
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1694700623
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_107
timestamp 1694700623
transform 1 0 13328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_139
timestamp 1694700623
transform 1 0 16912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_143
timestamp 1694700623
transform 1 0 17360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_145
timestamp 1694700623
transform 1 0 17584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_1671
timestamp 1694700623
transform 1 0 188496 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_1703
timestamp 1694700623
transform 1 0 192080 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1706
timestamp 1694700623
transform 1 0 192416 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1770
timestamp 1694700623
transform 1 0 199584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_1776
timestamp 1694700623
transform 1 0 200256 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1808
timestamp 1694700623
transform 1 0 203840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_1812
timestamp 1694700623
transform 1 0 204288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1694700623
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_12
timestamp 1694700623
transform 1 0 2688 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_44
timestamp 1694700623
transform 1 0 6272 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1694700623
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1694700623
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1694700623
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1694700623
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1694700623
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1671
timestamp 1694700623
transform 1 0 188496 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1735
timestamp 1694700623
transform 1 0 195664 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1741
timestamp 1694700623
transform 1 0 196336 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1805
timestamp 1694700623
transform 1 0 203504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_1811
timestamp 1694700623
transform 1 0 204176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_1813
timestamp 1694700623
transform 1 0 204400 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1694700623
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1694700623
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1694700623
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1694700623
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_107
timestamp 1694700623
transform 1 0 13328 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_139
timestamp 1694700623
transform 1 0 16912 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_143
timestamp 1694700623
transform 1 0 17360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_145
timestamp 1694700623
transform 1 0 17584 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_1671
timestamp 1694700623
transform 1 0 188496 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_1703
timestamp 1694700623
transform 1 0 192080 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1706
timestamp 1694700623
transform 1 0 192416 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1770
timestamp 1694700623
transform 1 0 199584 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_1776
timestamp 1694700623
transform 1 0 200256 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1808
timestamp 1694700623
transform 1 0 203840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_1812
timestamp 1694700623
transform 1 0 204288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1694700623
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1694700623
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1694700623
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1694700623
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1694700623
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1671
timestamp 1694700623
transform 1 0 188496 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1735
timestamp 1694700623
transform 1 0 195664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1741
timestamp 1694700623
transform 1 0 196336 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1805
timestamp 1694700623
transform 1 0 203504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_1811
timestamp 1694700623
transform 1 0 204176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_1813
timestamp 1694700623
transform 1 0 204400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1694700623
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1694700623
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1694700623
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1694700623
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1694700623
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_139
timestamp 1694700623
transform 1 0 16912 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_143
timestamp 1694700623
transform 1 0 17360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_145
timestamp 1694700623
transform 1 0 17584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_1671
timestamp 1694700623
transform 1 0 188496 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_1703
timestamp 1694700623
transform 1 0 192080 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1706
timestamp 1694700623
transform 1 0 192416 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1770
timestamp 1694700623
transform 1 0 199584 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_1776
timestamp 1694700623
transform 1 0 200256 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_1808
timestamp 1694700623
transform 1 0 203840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1694700623
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1694700623
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1694700623
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1694700623
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1694700623
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1671
timestamp 1694700623
transform 1 0 188496 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1735
timestamp 1694700623
transform 1 0 195664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1741
timestamp 1694700623
transform 1 0 196336 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1805
timestamp 1694700623
transform 1 0 203504 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_1811
timestamp 1694700623
transform 1 0 204176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_1813
timestamp 1694700623
transform 1 0 204400 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_6
timestamp 1694700623
transform 1 0 2016 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_22
timestamp 1694700623
transform 1 0 3808 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_30
timestamp 1694700623
transform 1 0 4704 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1694700623
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1694700623
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1694700623
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1694700623
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_139
timestamp 1694700623
transform 1 0 16912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_143
timestamp 1694700623
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_145
timestamp 1694700623
transform 1 0 17584 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_1671
timestamp 1694700623
transform 1 0 188496 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_1703
timestamp 1694700623
transform 1 0 192080 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1706
timestamp 1694700623
transform 1 0 192416 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1770
timestamp 1694700623
transform 1 0 199584 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_1776
timestamp 1694700623
transform 1 0 200256 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1808
timestamp 1694700623
transform 1 0 203840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_1812
timestamp 1694700623
transform 1 0 204288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1694700623
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1694700623
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1694700623
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1694700623
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1694700623
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1671
timestamp 1694700623
transform 1 0 188496 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1735
timestamp 1694700623
transform 1 0 195664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1741
timestamp 1694700623
transform 1 0 196336 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1805
timestamp 1694700623
transform 1 0 203504 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_1811
timestamp 1694700623
transform 1 0 204176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_1813
timestamp 1694700623
transform 1 0 204400 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1694700623
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1694700623
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1694700623
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1694700623
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1694700623
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_139
timestamp 1694700623
transform 1 0 16912 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_143
timestamp 1694700623
transform 1 0 17360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_145
timestamp 1694700623
transform 1 0 17584 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_1671
timestamp 1694700623
transform 1 0 188496 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_1703
timestamp 1694700623
transform 1 0 192080 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1706
timestamp 1694700623
transform 1 0 192416 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1770
timestamp 1694700623
transform 1 0 199584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_1776
timestamp 1694700623
transform 1 0 200256 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1808
timestamp 1694700623
transform 1 0 203840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_1812
timestamp 1694700623
transform 1 0 204288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1694700623
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1694700623
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1694700623
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1694700623
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_142
timestamp 1694700623
transform 1 0 17248 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1671
timestamp 1694700623
transform 1 0 188496 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1735
timestamp 1694700623
transform 1 0 195664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1741
timestamp 1694700623
transform 1 0 196336 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1805
timestamp 1694700623
transform 1 0 203504 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_1811
timestamp 1694700623
transform 1 0 204176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_1813
timestamp 1694700623
transform 1 0 204400 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_6
timestamp 1694700623
transform 1 0 2016 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_22
timestamp 1694700623
transform 1 0 3808 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_30
timestamp 1694700623
transform 1 0 4704 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1694700623
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1694700623
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1694700623
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1694700623
transform 1 0 13328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_139
timestamp 1694700623
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1694700623
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_145
timestamp 1694700623
transform 1 0 17584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_1671
timestamp 1694700623
transform 1 0 188496 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_1703
timestamp 1694700623
transform 1 0 192080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1706
timestamp 1694700623
transform 1 0 192416 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1770
timestamp 1694700623
transform 1 0 199584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_1776
timestamp 1694700623
transform 1 0 200256 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1808
timestamp 1694700623
transform 1 0 203840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_1812
timestamp 1694700623
transform 1 0 204288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1694700623
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1694700623
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1694700623
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1694700623
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1694700623
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1671
timestamp 1694700623
transform 1 0 188496 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1735
timestamp 1694700623
transform 1 0 195664 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1741
timestamp 1694700623
transform 1 0 196336 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1805
timestamp 1694700623
transform 1 0 203504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1811
timestamp 1694700623
transform 1 0 204176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_1813
timestamp 1694700623
transform 1 0 204400 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1694700623
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1694700623
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1694700623
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1694700623
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_107
timestamp 1694700623
transform 1 0 13328 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_139
timestamp 1694700623
transform 1 0 16912 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_143
timestamp 1694700623
transform 1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_145
timestamp 1694700623
transform 1 0 17584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_1671
timestamp 1694700623
transform 1 0 188496 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1703
timestamp 1694700623
transform 1 0 192080 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1706
timestamp 1694700623
transform 1 0 192416 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1770
timestamp 1694700623
transform 1 0 199584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_1776
timestamp 1694700623
transform 1 0 200256 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1808
timestamp 1694700623
transform 1 0 203840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1812
timestamp 1694700623
transform 1 0 204288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1694700623
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1694700623
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1694700623
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1694700623
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_142
timestamp 1694700623
transform 1 0 17248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1671
timestamp 1694700623
transform 1 0 188496 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1735
timestamp 1694700623
transform 1 0 195664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1741
timestamp 1694700623
transform 1 0 196336 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1805
timestamp 1694700623
transform 1 0 203504 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1811
timestamp 1694700623
transform 1 0 204176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_1813
timestamp 1694700623
transform 1 0 204400 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1694700623
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1694700623
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1694700623
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1694700623
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_107
timestamp 1694700623
transform 1 0 13328 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_139
timestamp 1694700623
transform 1 0 16912 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_143
timestamp 1694700623
transform 1 0 17360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_145
timestamp 1694700623
transform 1 0 17584 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_1671
timestamp 1694700623
transform 1 0 188496 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_1703
timestamp 1694700623
transform 1 0 192080 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1706
timestamp 1694700623
transform 1 0 192416 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1770
timestamp 1694700623
transform 1 0 199584 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_1776
timestamp 1694700623
transform 1 0 200256 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1808
timestamp 1694700623
transform 1 0 203840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_1812
timestamp 1694700623
transform 1 0 204288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_8
timestamp 1694700623
transform 1 0 2240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_12
timestamp 1694700623
transform 1 0 2688 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_44
timestamp 1694700623
transform 1 0 6272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_60
timestamp 1694700623
transform 1 0 8064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1694700623
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1694700623
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1694700623
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_142
timestamp 1694700623
transform 1 0 17248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1671
timestamp 1694700623
transform 1 0 188496 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1735
timestamp 1694700623
transform 1 0 195664 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1741
timestamp 1694700623
transform 1 0 196336 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1805
timestamp 1694700623
transform 1 0 203504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_1811
timestamp 1694700623
transform 1 0 204176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_1813
timestamp 1694700623
transform 1 0 204400 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1694700623
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1694700623
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1694700623
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1694700623
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_107
timestamp 1694700623
transform 1 0 13328 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_139
timestamp 1694700623
transform 1 0 16912 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_143
timestamp 1694700623
transform 1 0 17360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_145
timestamp 1694700623
transform 1 0 17584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_1671
timestamp 1694700623
transform 1 0 188496 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_1703
timestamp 1694700623
transform 1 0 192080 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1706
timestamp 1694700623
transform 1 0 192416 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1770
timestamp 1694700623
transform 1 0 199584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_1776
timestamp 1694700623
transform 1 0 200256 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1808
timestamp 1694700623
transform 1 0 203840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_1812
timestamp 1694700623
transform 1 0 204288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1694700623
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1694700623
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1694700623
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1694700623
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_142
timestamp 1694700623
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1671
timestamp 1694700623
transform 1 0 188496 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1735
timestamp 1694700623
transform 1 0 195664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1741
timestamp 1694700623
transform 1 0 196336 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1805
timestamp 1694700623
transform 1 0 203504 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_1811
timestamp 1694700623
transform 1 0 204176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_1813
timestamp 1694700623
transform 1 0 204400 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1694700623
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1694700623
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1694700623
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1694700623
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_107
timestamp 1694700623
transform 1 0 13328 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_139
timestamp 1694700623
transform 1 0 16912 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_143
timestamp 1694700623
transform 1 0 17360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_145
timestamp 1694700623
transform 1 0 17584 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_1671
timestamp 1694700623
transform 1 0 188496 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_1703
timestamp 1694700623
transform 1 0 192080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1706
timestamp 1694700623
transform 1 0 192416 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1770
timestamp 1694700623
transform 1 0 199584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_1776
timestamp 1694700623
transform 1 0 200256 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1808
timestamp 1694700623
transform 1 0 203840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_1812
timestamp 1694700623
transform 1 0 204288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1694700623
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1694700623
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1694700623
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_136
timestamp 1694700623
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1694700623
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1671
timestamp 1694700623
transform 1 0 188496 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1735
timestamp 1694700623
transform 1 0 195664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1741
timestamp 1694700623
transform 1 0 196336 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1805
timestamp 1694700623
transform 1 0 203504 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_1811
timestamp 1694700623
transform 1 0 204176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_1813
timestamp 1694700623
transform 1 0 204400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1694700623
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1694700623
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1694700623
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1694700623
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1694700623
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1694700623
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1694700623
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_139
timestamp 1694700623
transform 1 0 16912 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_143
timestamp 1694700623
transform 1 0 17360 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_1671
timestamp 1694700623
transform 1 0 188496 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_1703
timestamp 1694700623
transform 1 0 192080 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1706
timestamp 1694700623
transform 1 0 192416 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1770
timestamp 1694700623
transform 1 0 199584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_1776
timestamp 1694700623
transform 1 0 200256 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1808
timestamp 1694700623
transform 1 0 203840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_1812
timestamp 1694700623
transform 1 0 204288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1694700623
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1694700623
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1694700623
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1694700623
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_142
timestamp 1694700623
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1671
timestamp 1694700623
transform 1 0 188496 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1735
timestamp 1694700623
transform 1 0 195664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1741
timestamp 1694700623
transform 1 0 196336 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1805
timestamp 1694700623
transform 1 0 203504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_1811
timestamp 1694700623
transform 1 0 204176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_1813
timestamp 1694700623
transform 1 0 204400 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1694700623
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1694700623
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1694700623
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1694700623
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_107
timestamp 1694700623
transform 1 0 13328 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_139
timestamp 1694700623
transform 1 0 16912 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_143
timestamp 1694700623
transform 1 0 17360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_145
timestamp 1694700623
transform 1 0 17584 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_1671
timestamp 1694700623
transform 1 0 188496 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_1703
timestamp 1694700623
transform 1 0 192080 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1706
timestamp 1694700623
transform 1 0 192416 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1770
timestamp 1694700623
transform 1 0 199584 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_1776
timestamp 1694700623
transform 1 0 200256 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1808
timestamp 1694700623
transform 1 0 203840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_1812
timestamp 1694700623
transform 1 0 204288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1694700623
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1694700623
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1694700623
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1694700623
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1694700623
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_1671
timestamp 1694700623
transform 1 0 188496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1675
timestamp 1694700623
transform 1 0 188944 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1741
timestamp 1694700623
transform 1 0 196336 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1805
timestamp 1694700623
transform 1 0 203504 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_1811
timestamp 1694700623
transform 1 0 204176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_1813
timestamp 1694700623
transform 1 0 204400 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1694700623
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1694700623
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1694700623
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1694700623
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_107
timestamp 1694700623
transform 1 0 13328 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_139
timestamp 1694700623
transform 1 0 16912 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_143
timestamp 1694700623
transform 1 0 17360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_145
timestamp 1694700623
transform 1 0 17584 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_1671
timestamp 1694700623
transform 1 0 188496 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_1703
timestamp 1694700623
transform 1 0 192080 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1706
timestamp 1694700623
transform 1 0 192416 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1770
timestamp 1694700623
transform 1 0 199584 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_1776
timestamp 1694700623
transform 1 0 200256 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1808
timestamp 1694700623
transform 1 0 203840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_1812
timestamp 1694700623
transform 1 0 204288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_6
timestamp 1694700623
transform 1 0 2016 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1694700623
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1694700623
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_142
timestamp 1694700623
transform 1 0 17248 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1671
timestamp 1694700623
transform 1 0 188496 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1735
timestamp 1694700623
transform 1 0 195664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1741
timestamp 1694700623
transform 1 0 196336 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1805
timestamp 1694700623
transform 1 0 203504 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_1811
timestamp 1694700623
transform 1 0 204176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_1813
timestamp 1694700623
transform 1 0 204400 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1694700623
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1694700623
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1694700623
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1694700623
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_107
timestamp 1694700623
transform 1 0 13328 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_139
timestamp 1694700623
transform 1 0 16912 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_143
timestamp 1694700623
transform 1 0 17360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_145
timestamp 1694700623
transform 1 0 17584 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_1671
timestamp 1694700623
transform 1 0 188496 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_1703
timestamp 1694700623
transform 1 0 192080 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1706
timestamp 1694700623
transform 1 0 192416 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1770
timestamp 1694700623
transform 1 0 199584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_1776
timestamp 1694700623
transform 1 0 200256 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_1784
timestamp 1694700623
transform 1 0 201152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1694700623
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1694700623
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1694700623
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1694700623
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1694700623
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1671
timestamp 1694700623
transform 1 0 188496 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1735
timestamp 1694700623
transform 1 0 195664 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1741
timestamp 1694700623
transform 1 0 196336 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1805
timestamp 1694700623
transform 1 0 203504 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_1811
timestamp 1694700623
transform 1 0 204176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_1813
timestamp 1694700623
transform 1 0 204400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1694700623
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1694700623
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1694700623
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1694700623
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_107
timestamp 1694700623
transform 1 0 13328 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_139
timestamp 1694700623
transform 1 0 16912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_143
timestamp 1694700623
transform 1 0 17360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_145
timestamp 1694700623
transform 1 0 17584 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_1671
timestamp 1694700623
transform 1 0 188496 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_1703
timestamp 1694700623
transform 1 0 192080 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1706
timestamp 1694700623
transform 1 0 192416 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1770
timestamp 1694700623
transform 1 0 199584 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_1776
timestamp 1694700623
transform 1 0 200256 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1808
timestamp 1694700623
transform 1 0 203840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_1812
timestamp 1694700623
transform 1 0 204288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1694700623
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_6
timestamp 1694700623
transform 1 0 2016 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1694700623
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1694700623
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1694700623
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1671
timestamp 1694700623
transform 1 0 188496 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1735
timestamp 1694700623
transform 1 0 195664 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1741
timestamp 1694700623
transform 1 0 196336 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1805
timestamp 1694700623
transform 1 0 203504 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_1811
timestamp 1694700623
transform 1 0 204176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_1813
timestamp 1694700623
transform 1 0 204400 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_10
timestamp 1694700623
transform 1 0 2464 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_26
timestamp 1694700623
transform 1 0 4256 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1694700623
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1694700623
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1694700623
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_107
timestamp 1694700623
transform 1 0 13328 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_139
timestamp 1694700623
transform 1 0 16912 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_143
timestamp 1694700623
transform 1 0 17360 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_145
timestamp 1694700623
transform 1 0 17584 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_1671
timestamp 1694700623
transform 1 0 188496 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1703
timestamp 1694700623
transform 1 0 192080 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1706
timestamp 1694700623
transform 1 0 192416 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1770
timestamp 1694700623
transform 1 0 199584 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_1776
timestamp 1694700623
transform 1 0 200256 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1808
timestamp 1694700623
transform 1 0 203840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1812
timestamp 1694700623
transform 1 0 204288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1694700623
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1694700623
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1694700623
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1694700623
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_142
timestamp 1694700623
transform 1 0 17248 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1671
timestamp 1694700623
transform 1 0 188496 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1735
timestamp 1694700623
transform 1 0 195664 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1741
timestamp 1694700623
transform 1 0 196336 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1805
timestamp 1694700623
transform 1 0 203504 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1811
timestamp 1694700623
transform 1 0 204176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_1813
timestamp 1694700623
transform 1 0 204400 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1694700623
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1694700623
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1694700623
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1694700623
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_107
timestamp 1694700623
transform 1 0 13328 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_139
timestamp 1694700623
transform 1 0 16912 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_143
timestamp 1694700623
transform 1 0 17360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_145
timestamp 1694700623
transform 1 0 17584 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_1671
timestamp 1694700623
transform 1 0 188496 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1703
timestamp 1694700623
transform 1 0 192080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_1706
timestamp 1694700623
transform 1 0 192416 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1770
timestamp 1694700623
transform 1 0 199584 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_1776
timestamp 1694700623
transform 1 0 200256 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1808
timestamp 1694700623
transform 1 0 203840 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1812
timestamp 1694700623
transform 1 0 204288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1694700623
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1694700623
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1694700623
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1694700623
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_142
timestamp 1694700623
transform 1 0 17248 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1671
timestamp 1694700623
transform 1 0 188496 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1735
timestamp 1694700623
transform 1 0 195664 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_1741
timestamp 1694700623
transform 1 0 196336 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_1805
timestamp 1694700623
transform 1 0 203504 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_1811
timestamp 1694700623
transform 1 0 204176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_1813
timestamp 1694700623
transform 1 0 204400 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1694700623
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1694700623
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1694700623
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1694700623
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_107
timestamp 1694700623
transform 1 0 13328 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_139
timestamp 1694700623
transform 1 0 16912 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_143
timestamp 1694700623
transform 1 0 17360 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_145
timestamp 1694700623
transform 1 0 17584 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_1671
timestamp 1694700623
transform 1 0 188496 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_1703
timestamp 1694700623
transform 1 0 192080 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_1706
timestamp 1694700623
transform 1 0 192416 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1770
timestamp 1694700623
transform 1 0 199584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_1776
timestamp 1694700623
transform 1 0 200256 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_1808
timestamp 1694700623
transform 1 0 203840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_1812
timestamp 1694700623
transform 1 0 204288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_6
timestamp 1694700623
transform 1 0 2016 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1694700623
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1694700623
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_142
timestamp 1694700623
transform 1 0 17248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1671
timestamp 1694700623
transform 1 0 188496 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1735
timestamp 1694700623
transform 1 0 195664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_1741
timestamp 1694700623
transform 1 0 196336 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_1805
timestamp 1694700623
transform 1 0 203504 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_1811
timestamp 1694700623
transform 1 0 204176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_1813
timestamp 1694700623
transform 1 0 204400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1694700623
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1694700623
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1694700623
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1694700623
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_107
timestamp 1694700623
transform 1 0 13328 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_139
timestamp 1694700623
transform 1 0 16912 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_143
timestamp 1694700623
transform 1 0 17360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_145
timestamp 1694700623
transform 1 0 17584 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_1671
timestamp 1694700623
transform 1 0 188496 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_1703
timestamp 1694700623
transform 1 0 192080 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_1706
timestamp 1694700623
transform 1 0 192416 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1770
timestamp 1694700623
transform 1 0 199584 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_1776
timestamp 1694700623
transform 1 0 200256 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_1808
timestamp 1694700623
transform 1 0 203840 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_1812
timestamp 1694700623
transform 1 0 204288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1694700623
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1694700623
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1694700623
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1694700623
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_142
timestamp 1694700623
transform 1 0 17248 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1671
timestamp 1694700623
transform 1 0 188496 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_1735
timestamp 1694700623
transform 1 0 195664 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_1741
timestamp 1694700623
transform 1 0 196336 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_1811
timestamp 1694700623
transform 1 0 204176 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_1813
timestamp 1694700623
transform 1 0 204400 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1694700623
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1694700623
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1694700623
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1694700623
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_107
timestamp 1694700623
transform 1 0 13328 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_139
timestamp 1694700623
transform 1 0 16912 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_143
timestamp 1694700623
transform 1 0 17360 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_145
timestamp 1694700623
transform 1 0 17584 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_1671
timestamp 1694700623
transform 1 0 188496 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_1703
timestamp 1694700623
transform 1 0 192080 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_1706
timestamp 1694700623
transform 1 0 192416 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1770
timestamp 1694700623
transform 1 0 199584 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_1776
timestamp 1694700623
transform 1 0 200256 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_1808
timestamp 1694700623
transform 1 0 203840 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_1812
timestamp 1694700623
transform 1 0 204288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1694700623
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1694700623
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1694700623
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1694700623
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_142
timestamp 1694700623
transform 1 0 17248 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1671
timestamp 1694700623
transform 1 0 188496 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1735
timestamp 1694700623
transform 1 0 195664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_1741
timestamp 1694700623
transform 1 0 196336 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_1805
timestamp 1694700623
transform 1 0 203504 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_1811
timestamp 1694700623
transform 1 0 204176 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_1813
timestamp 1694700623
transform 1 0 204400 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_6
timestamp 1694700623
transform 1 0 2016 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_22
timestamp 1694700623
transform 1 0 3808 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_30
timestamp 1694700623
transform 1 0 4704 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1694700623
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1694700623
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1694700623
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_107
timestamp 1694700623
transform 1 0 13328 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_139
timestamp 1694700623
transform 1 0 16912 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_143
timestamp 1694700623
transform 1 0 17360 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_145
timestamp 1694700623
transform 1 0 17584 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_1671
timestamp 1694700623
transform 1 0 188496 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_1703
timestamp 1694700623
transform 1 0 192080 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_1706
timestamp 1694700623
transform 1 0 192416 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1770
timestamp 1694700623
transform 1 0 199584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_1776
timestamp 1694700623
transform 1 0 200256 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_1808
timestamp 1694700623
transform 1 0 203840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_1812
timestamp 1694700623
transform 1 0 204288 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1694700623
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1694700623
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1694700623
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1694700623
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_142
timestamp 1694700623
transform 1 0 17248 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1671
timestamp 1694700623
transform 1 0 188496 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1735
timestamp 1694700623
transform 1 0 195664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_1741
timestamp 1694700623
transform 1 0 196336 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_1805
timestamp 1694700623
transform 1 0 203504 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_1811
timestamp 1694700623
transform 1 0 204176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_1813
timestamp 1694700623
transform 1 0 204400 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1694700623
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1694700623
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1694700623
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1694700623
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_107
timestamp 1694700623
transform 1 0 13328 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_139
timestamp 1694700623
transform 1 0 16912 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_143
timestamp 1694700623
transform 1 0 17360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_145
timestamp 1694700623
transform 1 0 17584 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1671
timestamp 1694700623
transform 1 0 188496 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_1703
timestamp 1694700623
transform 1 0 192080 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_1706
timestamp 1694700623
transform 1 0 192416 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1770
timestamp 1694700623
transform 1 0 199584 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_1776
timestamp 1694700623
transform 1 0 200256 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_1808
timestamp 1694700623
transform 1 0 203840 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_1812
timestamp 1694700623
transform 1 0 204288 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_2
timestamp 1694700623
transform 1 0 1568 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_6
timestamp 1694700623
transform 1 0 2016 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1694700623
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1694700623
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_142
timestamp 1694700623
transform 1 0 17248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1671
timestamp 1694700623
transform 1 0 188496 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1735
timestamp 1694700623
transform 1 0 195664 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_1741
timestamp 1694700623
transform 1 0 196336 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_1805
timestamp 1694700623
transform 1 0 203504 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_1811
timestamp 1694700623
transform 1 0 204176 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_1813
timestamp 1694700623
transform 1 0 204400 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_10
timestamp 1694700623
transform 1 0 2464 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_26
timestamp 1694700623
transform 1 0 4256 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1694700623
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1694700623
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1694700623
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_107
timestamp 1694700623
transform 1 0 13328 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_139
timestamp 1694700623
transform 1 0 16912 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_143
timestamp 1694700623
transform 1 0 17360 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_145
timestamp 1694700623
transform 1 0 17584 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1671
timestamp 1694700623
transform 1 0 188496 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_1703
timestamp 1694700623
transform 1 0 192080 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_1706
timestamp 1694700623
transform 1 0 192416 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1770
timestamp 1694700623
transform 1 0 199584 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_1776
timestamp 1694700623
transform 1 0 200256 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_1808
timestamp 1694700623
transform 1 0 203840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_1812
timestamp 1694700623
transform 1 0 204288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_2
timestamp 1694700623
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_66
timestamp 1694700623
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1694700623
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1694700623
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_142
timestamp 1694700623
transform 1 0 17248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_1671
timestamp 1694700623
transform 1 0 188496 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1735
timestamp 1694700623
transform 1 0 195664 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_1741
timestamp 1694700623
transform 1 0 196336 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_1805
timestamp 1694700623
transform 1 0 203504 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_1811
timestamp 1694700623
transform 1 0 204176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_1813
timestamp 1694700623
transform 1 0 204400 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_2
timestamp 1694700623
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1694700623
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1694700623
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1694700623
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_107
timestamp 1694700623
transform 1 0 13328 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_139
timestamp 1694700623
transform 1 0 16912 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_143
timestamp 1694700623
transform 1 0 17360 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_145
timestamp 1694700623
transform 1 0 17584 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_1671
timestamp 1694700623
transform 1 0 188496 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_1703
timestamp 1694700623
transform 1 0 192080 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_1706
timestamp 1694700623
transform 1 0 192416 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_1770
timestamp 1694700623
transform 1 0 199584 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_1776
timestamp 1694700623
transform 1 0 200256 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_1808
timestamp 1694700623
transform 1 0 203840 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_1812
timestamp 1694700623
transform 1 0 204288 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_2
timestamp 1694700623
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1694700623
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1694700623
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1694700623
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_142
timestamp 1694700623
transform 1 0 17248 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_1671
timestamp 1694700623
transform 1 0 188496 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_1735
timestamp 1694700623
transform 1 0 195664 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_1741
timestamp 1694700623
transform 1 0 196336 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_1805
timestamp 1694700623
transform 1 0 203504 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_1811
timestamp 1694700623
transform 1 0 204176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_1813
timestamp 1694700623
transform 1 0 204400 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_2
timestamp 1694700623
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1694700623
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1694700623
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1694700623
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_107
timestamp 1694700623
transform 1 0 13328 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_139
timestamp 1694700623
transform 1 0 16912 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_143
timestamp 1694700623
transform 1 0 17360 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_145
timestamp 1694700623
transform 1 0 17584 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_1671
timestamp 1694700623
transform 1 0 188496 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_1703
timestamp 1694700623
transform 1 0 192080 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_1706
timestamp 1694700623
transform 1 0 192416 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_1770
timestamp 1694700623
transform 1 0 199584 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_1776
timestamp 1694700623
transform 1 0 200256 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_1808
timestamp 1694700623
transform 1 0 203840 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_1812
timestamp 1694700623
transform 1 0 204288 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_6
timestamp 1694700623
transform 1 0 2016 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1694700623
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1694700623
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_142
timestamp 1694700623
transform 1 0 17248 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_1671
timestamp 1694700623
transform 1 0 188496 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_1735
timestamp 1694700623
transform 1 0 195664 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_1741
timestamp 1694700623
transform 1 0 196336 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_1805
timestamp 1694700623
transform 1 0 203504 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_1811
timestamp 1694700623
transform 1 0 204176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_1813
timestamp 1694700623
transform 1 0 204400 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1694700623
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1694700623
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1694700623
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1694700623
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_107
timestamp 1694700623
transform 1 0 13328 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_139
timestamp 1694700623
transform 1 0 16912 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_143
timestamp 1694700623
transform 1 0 17360 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_145
timestamp 1694700623
transform 1 0 17584 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_1671
timestamp 1694700623
transform 1 0 188496 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_1703
timestamp 1694700623
transform 1 0 192080 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_1706
timestamp 1694700623
transform 1 0 192416 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_1770
timestamp 1694700623
transform 1 0 199584 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_1776
timestamp 1694700623
transform 1 0 200256 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_1808
timestamp 1694700623
transform 1 0 203840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_1812
timestamp 1694700623
transform 1 0 204288 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_2
timestamp 1694700623
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1694700623
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1694700623
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1694700623
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_142
timestamp 1694700623
transform 1 0 17248 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_1671
timestamp 1694700623
transform 1 0 188496 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_1735
timestamp 1694700623
transform 1 0 195664 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_1741
timestamp 1694700623
transform 1 0 196336 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_1805
timestamp 1694700623
transform 1 0 203504 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_1811
timestamp 1694700623
transform 1 0 204176 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_1813
timestamp 1694700623
transform 1 0 204400 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1694700623
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1694700623
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1694700623
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1694700623
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_107
timestamp 1694700623
transform 1 0 13328 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_139
timestamp 1694700623
transform 1 0 16912 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_143
timestamp 1694700623
transform 1 0 17360 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_145
timestamp 1694700623
transform 1 0 17584 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_1671
timestamp 1694700623
transform 1 0 188496 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_1703
timestamp 1694700623
transform 1 0 192080 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_1706
timestamp 1694700623
transform 1 0 192416 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_1770
timestamp 1694700623
transform 1 0 199584 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_1776
timestamp 1694700623
transform 1 0 200256 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_1808
timestamp 1694700623
transform 1 0 203840 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_1812
timestamp 1694700623
transform 1 0 204288 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_2
timestamp 1694700623
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_66
timestamp 1694700623
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1694700623
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1694700623
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_142
timestamp 1694700623
transform 1 0 17248 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_1671
timestamp 1694700623
transform 1 0 188496 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_1735
timestamp 1694700623
transform 1 0 195664 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_1741
timestamp 1694700623
transform 1 0 196336 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_1805
timestamp 1694700623
transform 1 0 203504 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_1811
timestamp 1694700623
transform 1 0 204176 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_1813
timestamp 1694700623
transform 1 0 204400 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_6
timestamp 1694700623
transform 1 0 2016 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_22
timestamp 1694700623
transform 1 0 3808 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_30
timestamp 1694700623
transform 1 0 4704 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1694700623
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1694700623
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1694700623
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_107
timestamp 1694700623
transform 1 0 13328 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_139
timestamp 1694700623
transform 1 0 16912 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_143
timestamp 1694700623
transform 1 0 17360 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_145
timestamp 1694700623
transform 1 0 17584 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_1671
timestamp 1694700623
transform 1 0 188496 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_1703
timestamp 1694700623
transform 1 0 192080 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_1706
timestamp 1694700623
transform 1 0 192416 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_1770
timestamp 1694700623
transform 1 0 199584 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_1776
timestamp 1694700623
transform 1 0 200256 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_1808
timestamp 1694700623
transform 1 0 203840 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_1812
timestamp 1694700623
transform 1 0 204288 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_2
timestamp 1694700623
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_66
timestamp 1694700623
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_72
timestamp 1694700623
transform 1 0 9408 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1694700623
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_142
timestamp 1694700623
transform 1 0 17248 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_1671
timestamp 1694700623
transform 1 0 188496 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_1735
timestamp 1694700623
transform 1 0 195664 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_1741
timestamp 1694700623
transform 1 0 196336 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_1805
timestamp 1694700623
transform 1 0 203504 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_1811
timestamp 1694700623
transform 1 0 204176 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_1813
timestamp 1694700623
transform 1 0 204400 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1694700623
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1694700623
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_37
timestamp 1694700623
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1694700623
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_107
timestamp 1694700623
transform 1 0 13328 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_139
timestamp 1694700623
transform 1 0 16912 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_143
timestamp 1694700623
transform 1 0 17360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_145
timestamp 1694700623
transform 1 0 17584 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_1671
timestamp 1694700623
transform 1 0 188496 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_1703
timestamp 1694700623
transform 1 0 192080 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_1706
timestamp 1694700623
transform 1 0 192416 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_1770
timestamp 1694700623
transform 1 0 199584 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_1776
timestamp 1694700623
transform 1 0 200256 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_1808
timestamp 1694700623
transform 1 0 203840 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_1812
timestamp 1694700623
transform 1 0 204288 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1694700623
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_66
timestamp 1694700623
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1694700623
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1694700623
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_142
timestamp 1694700623
transform 1 0 17248 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_1671
timestamp 1694700623
transform 1 0 188496 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_1735
timestamp 1694700623
transform 1 0 195664 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_1741
timestamp 1694700623
transform 1 0 196336 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_1805
timestamp 1694700623
transform 1 0 203504 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_1811
timestamp 1694700623
transform 1 0 204176 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_1813
timestamp 1694700623
transform 1 0 204400 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_2
timestamp 1694700623
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1694700623
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1694700623
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1694700623
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_107
timestamp 1694700623
transform 1 0 13328 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_139
timestamp 1694700623
transform 1 0 16912 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_143
timestamp 1694700623
transform 1 0 17360 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_145
timestamp 1694700623
transform 1 0 17584 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_1671
timestamp 1694700623
transform 1 0 188496 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_1703
timestamp 1694700623
transform 1 0 192080 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_1706
timestamp 1694700623
transform 1 0 192416 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_1770
timestamp 1694700623
transform 1 0 199584 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_1776
timestamp 1694700623
transform 1 0 200256 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_1808
timestamp 1694700623
transform 1 0 203840 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_1811
timestamp 1694700623
transform 1 0 204176 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_1813
timestamp 1694700623
transform 1 0 204400 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_8
timestamp 1694700623
transform 1 0 2240 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_12
timestamp 1694700623
transform 1 0 2688 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_44
timestamp 1694700623
transform 1 0 6272 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_60
timestamp 1694700623
transform 1 0 8064 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_68
timestamp 1694700623
transform 1 0 8960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_72
timestamp 1694700623
transform 1 0 9408 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_136
timestamp 1694700623
transform 1 0 16576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_142
timestamp 1694700623
transform 1 0 17248 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_1671
timestamp 1694700623
transform 1 0 188496 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_1735
timestamp 1694700623
transform 1 0 195664 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_1741
timestamp 1694700623
transform 1 0 196336 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_1773
timestamp 1694700623
transform 1 0 199920 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_1781
timestamp 1694700623
transform 1 0 200816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_1811
timestamp 1694700623
transform 1 0 204176 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_1813
timestamp 1694700623
transform 1 0 204400 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_2
timestamp 1694700623
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1694700623
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1694700623
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1694700623
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_107
timestamp 1694700623
transform 1 0 13328 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_139
timestamp 1694700623
transform 1 0 16912 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_143
timestamp 1694700623
transform 1 0 17360 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_145
timestamp 1694700623
transform 1 0 17584 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_1671
timestamp 1694700623
transform 1 0 188496 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_1703
timestamp 1694700623
transform 1 0 192080 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_1706
timestamp 1694700623
transform 1 0 192416 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_1770
timestamp 1694700623
transform 1 0 199584 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_1776
timestamp 1694700623
transform 1 0 200256 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_1808
timestamp 1694700623
transform 1 0 203840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_1812
timestamp 1694700623
transform 1 0 204288 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_2
timestamp 1694700623
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_66
timestamp 1694700623
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1694700623
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1694700623
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_142
timestamp 1694700623
transform 1 0 17248 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_1671
timestamp 1694700623
transform 1 0 188496 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_1735
timestamp 1694700623
transform 1 0 195664 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_1741
timestamp 1694700623
transform 1 0 196336 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_1805
timestamp 1694700623
transform 1 0 203504 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_1811
timestamp 1694700623
transform 1 0 204176 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_1813
timestamp 1694700623
transform 1 0 204400 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1694700623
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1694700623
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1694700623
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1694700623
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_107
timestamp 1694700623
transform 1 0 13328 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_139
timestamp 1694700623
transform 1 0 16912 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_143
timestamp 1694700623
transform 1 0 17360 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_145
timestamp 1694700623
transform 1 0 17584 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_1671
timestamp 1694700623
transform 1 0 188496 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_1703
timestamp 1694700623
transform 1 0 192080 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_1706
timestamp 1694700623
transform 1 0 192416 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_1770
timestamp 1694700623
transform 1 0 199584 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_1776
timestamp 1694700623
transform 1 0 200256 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_1808
timestamp 1694700623
transform 1 0 203840 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_1812
timestamp 1694700623
transform 1 0 204288 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_2
timestamp 1694700623
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_66
timestamp 1694700623
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1694700623
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1694700623
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_142
timestamp 1694700623
transform 1 0 17248 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_1671
timestamp 1694700623
transform 1 0 188496 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_1735
timestamp 1694700623
transform 1 0 195664 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_1741
timestamp 1694700623
transform 1 0 196336 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_1805
timestamp 1694700623
transform 1 0 203504 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_1811
timestamp 1694700623
transform 1 0 204176 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_1813
timestamp 1694700623
transform 1 0 204400 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_6
timestamp 1694700623
transform 1 0 2016 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_22
timestamp 1694700623
transform 1 0 3808 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_30
timestamp 1694700623
transform 1 0 4704 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1694700623
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1694700623
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1694700623
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_107
timestamp 1694700623
transform 1 0 13328 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_139
timestamp 1694700623
transform 1 0 16912 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_143
timestamp 1694700623
transform 1 0 17360 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_145
timestamp 1694700623
transform 1 0 17584 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_1671
timestamp 1694700623
transform 1 0 188496 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_1703
timestamp 1694700623
transform 1 0 192080 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_1706
timestamp 1694700623
transform 1 0 192416 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_1770
timestamp 1694700623
transform 1 0 199584 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_1776
timestamp 1694700623
transform 1 0 200256 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_1808
timestamp 1694700623
transform 1 0 203840 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_1812
timestamp 1694700623
transform 1 0 204288 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1694700623
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1694700623
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1694700623
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1694700623
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_142
timestamp 1694700623
transform 1 0 17248 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_1671
timestamp 1694700623
transform 1 0 188496 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_1735
timestamp 1694700623
transform 1 0 195664 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_1741
timestamp 1694700623
transform 1 0 196336 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_1805
timestamp 1694700623
transform 1 0 203504 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_1811
timestamp 1694700623
transform 1 0 204176 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_1813
timestamp 1694700623
transform 1 0 204400 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1694700623
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1694700623
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1694700623
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1694700623
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_107
timestamp 1694700623
transform 1 0 13328 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_139
timestamp 1694700623
transform 1 0 16912 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_143
timestamp 1694700623
transform 1 0 17360 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_145
timestamp 1694700623
transform 1 0 17584 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_1671
timestamp 1694700623
transform 1 0 188496 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_1703
timestamp 1694700623
transform 1 0 192080 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_1706
timestamp 1694700623
transform 1 0 192416 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_1770
timestamp 1694700623
transform 1 0 199584 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_1776
timestamp 1694700623
transform 1 0 200256 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_1808
timestamp 1694700623
transform 1 0 203840 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_1812
timestamp 1694700623
transform 1 0 204288 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_2
timestamp 1694700623
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1694700623
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_72
timestamp 1694700623
transform 1 0 9408 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_136
timestamp 1694700623
transform 1 0 16576 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_142
timestamp 1694700623
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_1671
timestamp 1694700623
transform 1 0 188496 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_1735
timestamp 1694700623
transform 1 0 195664 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_1741
timestamp 1694700623
transform 1 0 196336 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_1805
timestamp 1694700623
transform 1 0 203504 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_1811
timestamp 1694700623
transform 1 0 204176 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_1813
timestamp 1694700623
transform 1 0 204400 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1694700623
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1694700623
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_37
timestamp 1694700623
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1694700623
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_107
timestamp 1694700623
transform 1 0 13328 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_139
timestamp 1694700623
transform 1 0 16912 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_143
timestamp 1694700623
transform 1 0 17360 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_145
timestamp 1694700623
transform 1 0 17584 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_1671
timestamp 1694700623
transform 1 0 188496 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_1703
timestamp 1694700623
transform 1 0 192080 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_1706
timestamp 1694700623
transform 1 0 192416 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_1770
timestamp 1694700623
transform 1 0 199584 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_1776
timestamp 1694700623
transform 1 0 200256 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_1808
timestamp 1694700623
transform 1 0 203840 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_1812
timestamp 1694700623
transform 1 0 204288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_6
timestamp 1694700623
transform 1 0 2016 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_72
timestamp 1694700623
transform 1 0 9408 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_136
timestamp 1694700623
transform 1 0 16576 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_142
timestamp 1694700623
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_1671
timestamp 1694700623
transform 1 0 188496 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_1735
timestamp 1694700623
transform 1 0 195664 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_1741
timestamp 1694700623
transform 1 0 196336 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_1805
timestamp 1694700623
transform 1 0 203504 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_1811
timestamp 1694700623
transform 1 0 204176 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_1813
timestamp 1694700623
transform 1 0 204400 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1694700623
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1694700623
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_37
timestamp 1694700623
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_101
timestamp 1694700623
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_107
timestamp 1694700623
transform 1 0 13328 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_139
timestamp 1694700623
transform 1 0 16912 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_143
timestamp 1694700623
transform 1 0 17360 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_1671
timestamp 1694700623
transform 1 0 188496 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_1703
timestamp 1694700623
transform 1 0 192080 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_1706
timestamp 1694700623
transform 1 0 192416 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_1770
timestamp 1694700623
transform 1 0 199584 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_1776
timestamp 1694700623
transform 1 0 200256 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_1808
timestamp 1694700623
transform 1 0 203840 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_2
timestamp 1694700623
transform 1 0 1568 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_66
timestamp 1694700623
transform 1 0 8736 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_72
timestamp 1694700623
transform 1 0 9408 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_136
timestamp 1694700623
transform 1 0 16576 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_142
timestamp 1694700623
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_1671
timestamp 1694700623
transform 1 0 188496 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_1735
timestamp 1694700623
transform 1 0 195664 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_1741
timestamp 1694700623
transform 1 0 196336 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_1805
timestamp 1694700623
transform 1 0 203504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_1811
timestamp 1694700623
transform 1 0 204176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_1813
timestamp 1694700623
transform 1 0 204400 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_2
timestamp 1694700623
transform 1 0 1568 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_34
timestamp 1694700623
transform 1 0 5152 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_37
timestamp 1694700623
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_101
timestamp 1694700623
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_107
timestamp 1694700623
transform 1 0 13328 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_139
timestamp 1694700623
transform 1 0 16912 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_143
timestamp 1694700623
transform 1 0 17360 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_145
timestamp 1694700623
transform 1 0 17584 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_1671
timestamp 1694700623
transform 1 0 188496 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_1703
timestamp 1694700623
transform 1 0 192080 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_1706
timestamp 1694700623
transform 1 0 192416 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_1770
timestamp 1694700623
transform 1 0 199584 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_1776
timestamp 1694700623
transform 1 0 200256 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_1808
timestamp 1694700623
transform 1 0 203840 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_1812
timestamp 1694700623
transform 1 0 204288 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_2
timestamp 1694700623
transform 1 0 1568 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_66
timestamp 1694700623
transform 1 0 8736 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_72
timestamp 1694700623
transform 1 0 9408 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_136
timestamp 1694700623
transform 1 0 16576 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_142
timestamp 1694700623
transform 1 0 17248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_1671
timestamp 1694700623
transform 1 0 188496 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_1735
timestamp 1694700623
transform 1 0 195664 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_1741
timestamp 1694700623
transform 1 0 196336 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_1805
timestamp 1694700623
transform 1 0 203504 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_1811
timestamp 1694700623
transform 1 0 204176 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_1813
timestamp 1694700623
transform 1 0 204400 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_8
timestamp 1694700623
transform 1 0 2240 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_12
timestamp 1694700623
transform 1 0 2688 0 1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_28
timestamp 1694700623
transform 1 0 4480 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_32
timestamp 1694700623
transform 1 0 4928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_34
timestamp 1694700623
transform 1 0 5152 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_37
timestamp 1694700623
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_101
timestamp 1694700623
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_107
timestamp 1694700623
transform 1 0 13328 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_139
timestamp 1694700623
transform 1 0 16912 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_143
timestamp 1694700623
transform 1 0 17360 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_1671
timestamp 1694700623
transform 1 0 188496 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_1703
timestamp 1694700623
transform 1 0 192080 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_1706
timestamp 1694700623
transform 1 0 192416 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_1770
timestamp 1694700623
transform 1 0 199584 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_1776
timestamp 1694700623
transform 1 0 200256 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_1808
timestamp 1694700623
transform 1 0 203840 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_1812
timestamp 1694700623
transform 1 0 204288 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_2
timestamp 1694700623
transform 1 0 1568 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_66
timestamp 1694700623
transform 1 0 8736 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_72
timestamp 1694700623
transform 1 0 9408 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_136
timestamp 1694700623
transform 1 0 16576 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_142
timestamp 1694700623
transform 1 0 17248 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_1671
timestamp 1694700623
transform 1 0 188496 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_1735
timestamp 1694700623
transform 1 0 195664 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_1741
timestamp 1694700623
transform 1 0 196336 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_1805
timestamp 1694700623
transform 1 0 203504 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_1811
timestamp 1694700623
transform 1 0 204176 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_1813
timestamp 1694700623
transform 1 0 204400 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_2
timestamp 1694700623
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_34
timestamp 1694700623
transform 1 0 5152 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_37
timestamp 1694700623
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_101
timestamp 1694700623
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_107
timestamp 1694700623
transform 1 0 13328 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_139
timestamp 1694700623
transform 1 0 16912 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_143
timestamp 1694700623
transform 1 0 17360 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_145
timestamp 1694700623
transform 1 0 17584 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_1671
timestamp 1694700623
transform 1 0 188496 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_1703
timestamp 1694700623
transform 1 0 192080 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_1706
timestamp 1694700623
transform 1 0 192416 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_1770
timestamp 1694700623
transform 1 0 199584 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_1776
timestamp 1694700623
transform 1 0 200256 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_1808
timestamp 1694700623
transform 1 0 203840 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_1812
timestamp 1694700623
transform 1 0 204288 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_2
timestamp 1694700623
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_66
timestamp 1694700623
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_72
timestamp 1694700623
transform 1 0 9408 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_136
timestamp 1694700623
transform 1 0 16576 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_142
timestamp 1694700623
transform 1 0 17248 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_1671
timestamp 1694700623
transform 1 0 188496 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_1735
timestamp 1694700623
transform 1 0 195664 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_1741
timestamp 1694700623
transform 1 0 196336 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_1805
timestamp 1694700623
transform 1 0 203504 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_1811
timestamp 1694700623
transform 1 0 204176 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_1813
timestamp 1694700623
transform 1 0 204400 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_6
timestamp 1694700623
transform 1 0 2016 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_22
timestamp 1694700623
transform 1 0 3808 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_30
timestamp 1694700623
transform 1 0 4704 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_34
timestamp 1694700623
transform 1 0 5152 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_37
timestamp 1694700623
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_101
timestamp 1694700623
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_107
timestamp 1694700623
transform 1 0 13328 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_139
timestamp 1694700623
transform 1 0 16912 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_143
timestamp 1694700623
transform 1 0 17360 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_145
timestamp 1694700623
transform 1 0 17584 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_1671
timestamp 1694700623
transform 1 0 188496 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_1703
timestamp 1694700623
transform 1 0 192080 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_1706
timestamp 1694700623
transform 1 0 192416 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_1770
timestamp 1694700623
transform 1 0 199584 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_1776
timestamp 1694700623
transform 1 0 200256 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_1808
timestamp 1694700623
transform 1 0 203840 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_1812
timestamp 1694700623
transform 1 0 204288 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_2
timestamp 1694700623
transform 1 0 1568 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_66
timestamp 1694700623
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_72
timestamp 1694700623
transform 1 0 9408 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_136
timestamp 1694700623
transform 1 0 16576 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_142
timestamp 1694700623
transform 1 0 17248 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_1671
timestamp 1694700623
transform 1 0 188496 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_1735
timestamp 1694700623
transform 1 0 195664 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_1741
timestamp 1694700623
transform 1 0 196336 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_1805
timestamp 1694700623
transform 1 0 203504 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_1811
timestamp 1694700623
transform 1 0 204176 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_1813
timestamp 1694700623
transform 1 0 204400 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_2
timestamp 1694700623
transform 1 0 1568 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_34
timestamp 1694700623
transform 1 0 5152 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_37
timestamp 1694700623
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_101
timestamp 1694700623
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_107
timestamp 1694700623
transform 1 0 13328 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_139
timestamp 1694700623
transform 1 0 16912 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_143
timestamp 1694700623
transform 1 0 17360 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_145
timestamp 1694700623
transform 1 0 17584 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_1671
timestamp 1694700623
transform 1 0 188496 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_1703
timestamp 1694700623
transform 1 0 192080 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_1706
timestamp 1694700623
transform 1 0 192416 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_1770
timestamp 1694700623
transform 1 0 199584 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_1776
timestamp 1694700623
transform 1 0 200256 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_1808
timestamp 1694700623
transform 1 0 203840 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_1812
timestamp 1694700623
transform 1 0 204288 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_2
timestamp 1694700623
transform 1 0 1568 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_66
timestamp 1694700623
transform 1 0 8736 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_72
timestamp 1694700623
transform 1 0 9408 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_136
timestamp 1694700623
transform 1 0 16576 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_142
timestamp 1694700623
transform 1 0 17248 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_1671
timestamp 1694700623
transform 1 0 188496 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_1735
timestamp 1694700623
transform 1 0 195664 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_1741
timestamp 1694700623
transform 1 0 196336 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_1805
timestamp 1694700623
transform 1 0 203504 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_1811
timestamp 1694700623
transform 1 0 204176 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_1813
timestamp 1694700623
transform 1 0 204400 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_2
timestamp 1694700623
transform 1 0 1568 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_34
timestamp 1694700623
transform 1 0 5152 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_37
timestamp 1694700623
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_101
timestamp 1694700623
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_107
timestamp 1694700623
transform 1 0 13328 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_139
timestamp 1694700623
transform 1 0 16912 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_143
timestamp 1694700623
transform 1 0 17360 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_145
timestamp 1694700623
transform 1 0 17584 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_1671
timestamp 1694700623
transform 1 0 188496 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_1703
timestamp 1694700623
transform 1 0 192080 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_1706
timestamp 1694700623
transform 1 0 192416 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_1770
timestamp 1694700623
transform 1 0 199584 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_1776
timestamp 1694700623
transform 1 0 200256 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_1808
timestamp 1694700623
transform 1 0 203840 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_1812
timestamp 1694700623
transform 1 0 204288 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_6
timestamp 1694700623
transform 1 0 2016 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_72
timestamp 1694700623
transform 1 0 9408 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_136
timestamp 1694700623
transform 1 0 16576 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_142
timestamp 1694700623
transform 1 0 17248 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_1671
timestamp 1694700623
transform 1 0 188496 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_1735
timestamp 1694700623
transform 1 0 195664 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_1741
timestamp 1694700623
transform 1 0 196336 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_1805
timestamp 1694700623
transform 1 0 203504 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_1811
timestamp 1694700623
transform 1 0 204176 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_1813
timestamp 1694700623
transform 1 0 204400 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_106_2
timestamp 1694700623
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_34
timestamp 1694700623
transform 1 0 5152 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_37
timestamp 1694700623
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_101
timestamp 1694700623
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_106_107
timestamp 1694700623
transform 1 0 13328 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_139
timestamp 1694700623
transform 1 0 16912 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_143
timestamp 1694700623
transform 1 0 17360 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_145
timestamp 1694700623
transform 1 0 17584 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_106_1671
timestamp 1694700623
transform 1 0 188496 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_1703
timestamp 1694700623
transform 1 0 192080 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_1706
timestamp 1694700623
transform 1 0 192416 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_1770
timestamp 1694700623
transform 1 0 199584 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_106_1776
timestamp 1694700623
transform 1 0 200256 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_1808
timestamp 1694700623
transform 1 0 203840 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_1812
timestamp 1694700623
transform 1 0 204288 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_2
timestamp 1694700623
transform 1 0 1568 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_66
timestamp 1694700623
transform 1 0 8736 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_72
timestamp 1694700623
transform 1 0 9408 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_136
timestamp 1694700623
transform 1 0 16576 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_142
timestamp 1694700623
transform 1 0 17248 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_1671
timestamp 1694700623
transform 1 0 188496 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_1735
timestamp 1694700623
transform 1 0 195664 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_1741
timestamp 1694700623
transform 1 0 196336 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_1805
timestamp 1694700623
transform 1 0 203504 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_1811
timestamp 1694700623
transform 1 0 204176 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_1813
timestamp 1694700623
transform 1 0 204400 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_2
timestamp 1694700623
transform 1 0 1568 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_34
timestamp 1694700623
transform 1 0 5152 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_37
timestamp 1694700623
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_101
timestamp 1694700623
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_107
timestamp 1694700623
transform 1 0 13328 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_139
timestamp 1694700623
transform 1 0 16912 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_143
timestamp 1694700623
transform 1 0 17360 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_145
timestamp 1694700623
transform 1 0 17584 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_1671
timestamp 1694700623
transform 1 0 188496 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_1703
timestamp 1694700623
transform 1 0 192080 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_1706
timestamp 1694700623
transform 1 0 192416 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_1770
timestamp 1694700623
transform 1 0 199584 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_1776
timestamp 1694700623
transform 1 0 200256 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_1808
timestamp 1694700623
transform 1 0 203840 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_1812
timestamp 1694700623
transform 1 0 204288 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_2
timestamp 1694700623
transform 1 0 1568 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_66
timestamp 1694700623
transform 1 0 8736 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_72
timestamp 1694700623
transform 1 0 9408 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_136
timestamp 1694700623
transform 1 0 16576 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_142
timestamp 1694700623
transform 1 0 17248 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_1671
timestamp 1694700623
transform 1 0 188496 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_1735
timestamp 1694700623
transform 1 0 195664 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_1741
timestamp 1694700623
transform 1 0 196336 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_1805
timestamp 1694700623
transform 1 0 203504 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_1811
timestamp 1694700623
transform 1 0 204176 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_1813
timestamp 1694700623
transform 1 0 204400 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_8
timestamp 1694700623
transform 1 0 2240 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_110_12
timestamp 1694700623
transform 1 0 2688 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_28
timestamp 1694700623
transform 1 0 4480 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_32
timestamp 1694700623
transform 1 0 4928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_34
timestamp 1694700623
transform 1 0 5152 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_37
timestamp 1694700623
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_101
timestamp 1694700623
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_110_107
timestamp 1694700623
transform 1 0 13328 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_139
timestamp 1694700623
transform 1 0 16912 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_143
timestamp 1694700623
transform 1 0 17360 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_145
timestamp 1694700623
transform 1 0 17584 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_110_1671
timestamp 1694700623
transform 1 0 188496 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_1703
timestamp 1694700623
transform 1 0 192080 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_1706
timestamp 1694700623
transform 1 0 192416 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_1770
timestamp 1694700623
transform 1 0 199584 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_110_1776
timestamp 1694700623
transform 1 0 200256 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_1808
timestamp 1694700623
transform 1 0 203840 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_1812
timestamp 1694700623
transform 1 0 204288 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_2
timestamp 1694700623
transform 1 0 1568 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_66
timestamp 1694700623
transform 1 0 8736 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_72
timestamp 1694700623
transform 1 0 9408 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_136
timestamp 1694700623
transform 1 0 16576 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_142
timestamp 1694700623
transform 1 0 17248 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_1671
timestamp 1694700623
transform 1 0 188496 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_1735
timestamp 1694700623
transform 1 0 195664 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_1741
timestamp 1694700623
transform 1 0 196336 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_1805
timestamp 1694700623
transform 1 0 203504 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_1811
timestamp 1694700623
transform 1 0 204176 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_1813
timestamp 1694700623
transform 1 0 204400 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_2
timestamp 1694700623
transform 1 0 1568 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_34
timestamp 1694700623
transform 1 0 5152 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_37
timestamp 1694700623
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_101
timestamp 1694700623
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_107
timestamp 1694700623
transform 1 0 13328 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_139
timestamp 1694700623
transform 1 0 16912 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_143
timestamp 1694700623
transform 1 0 17360 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_145
timestamp 1694700623
transform 1 0 17584 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_1671
timestamp 1694700623
transform 1 0 188496 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_1703
timestamp 1694700623
transform 1 0 192080 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_1706
timestamp 1694700623
transform 1 0 192416 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_1770
timestamp 1694700623
transform 1 0 199584 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_1776
timestamp 1694700623
transform 1 0 200256 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_1808
timestamp 1694700623
transform 1 0 203840 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_1812
timestamp 1694700623
transform 1 0 204288 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_2
timestamp 1694700623
transform 1 0 1568 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_66
timestamp 1694700623
transform 1 0 8736 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_72
timestamp 1694700623
transform 1 0 9408 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_136
timestamp 1694700623
transform 1 0 16576 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_142
timestamp 1694700623
transform 1 0 17248 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_1671
timestamp 1694700623
transform 1 0 188496 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_1735
timestamp 1694700623
transform 1 0 195664 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_1741
timestamp 1694700623
transform 1 0 196336 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_1805
timestamp 1694700623
transform 1 0 203504 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_1811
timestamp 1694700623
transform 1 0 204176 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_1813
timestamp 1694700623
transform 1 0 204400 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_2
timestamp 1694700623
transform 1 0 1568 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_34
timestamp 1694700623
transform 1 0 5152 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_37
timestamp 1694700623
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_101
timestamp 1694700623
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_107
timestamp 1694700623
transform 1 0 13328 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_139
timestamp 1694700623
transform 1 0 16912 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_143
timestamp 1694700623
transform 1 0 17360 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_145
timestamp 1694700623
transform 1 0 17584 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_1671
timestamp 1694700623
transform 1 0 188496 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_1703
timestamp 1694700623
transform 1 0 192080 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_1706
timestamp 1694700623
transform 1 0 192416 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_1770
timestamp 1694700623
transform 1 0 199584 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_1776
timestamp 1694700623
transform 1 0 200256 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_1808
timestamp 1694700623
transform 1 0 203840 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_1811
timestamp 1694700623
transform 1 0 204176 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_1813
timestamp 1694700623
transform 1 0 204400 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_6
timestamp 1694700623
transform 1 0 2016 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_72
timestamp 1694700623
transform 1 0 9408 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_136
timestamp 1694700623
transform 1 0 16576 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_142
timestamp 1694700623
transform 1 0 17248 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_1671
timestamp 1694700623
transform 1 0 188496 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_1735
timestamp 1694700623
transform 1 0 195664 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_115_1741
timestamp 1694700623
transform 1 0 196336 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_1773
timestamp 1694700623
transform 1 0 199920 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_1781
timestamp 1694700623
transform 1 0 200816 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_1811
timestamp 1694700623
transform 1 0 204176 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_1813
timestamp 1694700623
transform 1 0 204400 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_116_2
timestamp 1694700623
transform 1 0 1568 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_34
timestamp 1694700623
transform 1 0 5152 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_37
timestamp 1694700623
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_101
timestamp 1694700623
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_116_107
timestamp 1694700623
transform 1 0 13328 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_139
timestamp 1694700623
transform 1 0 16912 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_143
timestamp 1694700623
transform 1 0 17360 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_145
timestamp 1694700623
transform 1 0 17584 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_116_1671
timestamp 1694700623
transform 1 0 188496 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_1703
timestamp 1694700623
transform 1 0 192080 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_1706
timestamp 1694700623
transform 1 0 192416 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_1770
timestamp 1694700623
transform 1 0 199584 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_116_1776
timestamp 1694700623
transform 1 0 200256 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_1808
timestamp 1694700623
transform 1 0 203840 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_1812
timestamp 1694700623
transform 1 0 204288 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_2
timestamp 1694700623
transform 1 0 1568 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_66
timestamp 1694700623
transform 1 0 8736 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_72
timestamp 1694700623
transform 1 0 9408 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_136
timestamp 1694700623
transform 1 0 16576 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_142
timestamp 1694700623
transform 1 0 17248 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_1671
timestamp 1694700623
transform 1 0 188496 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_1735
timestamp 1694700623
transform 1 0 195664 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_1741
timestamp 1694700623
transform 1 0 196336 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_1805
timestamp 1694700623
transform 1 0 203504 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_1811
timestamp 1694700623
transform 1 0 204176 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_1813
timestamp 1694700623
transform 1 0 204400 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_2
timestamp 1694700623
transform 1 0 1568 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_34
timestamp 1694700623
transform 1 0 5152 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_118_37
timestamp 1694700623
transform 1 0 5488 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_101
timestamp 1694700623
transform 1 0 12656 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_107
timestamp 1694700623
transform 1 0 13328 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_139
timestamp 1694700623
transform 1 0 16912 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_143
timestamp 1694700623
transform 1 0 17360 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_145
timestamp 1694700623
transform 1 0 17584 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_1671
timestamp 1694700623
transform 1 0 188496 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_1703
timestamp 1694700623
transform 1 0 192080 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_118_1706
timestamp 1694700623
transform 1 0 192416 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_1770
timestamp 1694700623
transform 1 0 199584 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_1776
timestamp 1694700623
transform 1 0 200256 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_1808
timestamp 1694700623
transform 1 0 203840 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_1812
timestamp 1694700623
transform 1 0 204288 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_119_2
timestamp 1694700623
transform 1 0 1568 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_66
timestamp 1694700623
transform 1 0 8736 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_119_72
timestamp 1694700623
transform 1 0 9408 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_136
timestamp 1694700623
transform 1 0 16576 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_142
timestamp 1694700623
transform 1 0 17248 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_119_1671
timestamp 1694700623
transform 1 0 188496 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_1735
timestamp 1694700623
transform 1 0 195664 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_119_1741
timestamp 1694700623
transform 1 0 196336 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_1805
timestamp 1694700623
transform 1 0 203504 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_1811
timestamp 1694700623
transform 1 0 204176 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_1813
timestamp 1694700623
transform 1 0 204400 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_120_6
timestamp 1694700623
transform 1 0 2016 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_22
timestamp 1694700623
transform 1 0 3808 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_30
timestamp 1694700623
transform 1 0 4704 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_34
timestamp 1694700623
transform 1 0 5152 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_120_37
timestamp 1694700623
transform 1 0 5488 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_101
timestamp 1694700623
transform 1 0 12656 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_120_107
timestamp 1694700623
transform 1 0 13328 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_139
timestamp 1694700623
transform 1 0 16912 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_143
timestamp 1694700623
transform 1 0 17360 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_145
timestamp 1694700623
transform 1 0 17584 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_120_1671
timestamp 1694700623
transform 1 0 188496 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_1703
timestamp 1694700623
transform 1 0 192080 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_120_1706
timestamp 1694700623
transform 1 0 192416 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_1770
timestamp 1694700623
transform 1 0 199584 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_120_1776
timestamp 1694700623
transform 1 0 200256 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_1808
timestamp 1694700623
transform 1 0 203840 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_1812
timestamp 1694700623
transform 1 0 204288 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_121_2
timestamp 1694700623
transform 1 0 1568 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_66
timestamp 1694700623
transform 1 0 8736 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_121_72
timestamp 1694700623
transform 1 0 9408 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_136
timestamp 1694700623
transform 1 0 16576 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_142
timestamp 1694700623
transform 1 0 17248 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_121_1671
timestamp 1694700623
transform 1 0 188496 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_1735
timestamp 1694700623
transform 1 0 195664 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_121_1741
timestamp 1694700623
transform 1 0 196336 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_1805
timestamp 1694700623
transform 1 0 203504 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_1811
timestamp 1694700623
transform 1 0 204176 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_1813
timestamp 1694700623
transform 1 0 204400 0 -1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_2
timestamp 1694700623
transform 1 0 1568 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_34
timestamp 1694700623
transform 1 0 5152 0 1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_122_37
timestamp 1694700623
transform 1 0 5488 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_101
timestamp 1694700623
transform 1 0 12656 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_107
timestamp 1694700623
transform 1 0 13328 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_139
timestamp 1694700623
transform 1 0 16912 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_143
timestamp 1694700623
transform 1 0 17360 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_145
timestamp 1694700623
transform 1 0 17584 0 1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_1671
timestamp 1694700623
transform 1 0 188496 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_1703
timestamp 1694700623
transform 1 0 192080 0 1 98784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_122_1706
timestamp 1694700623
transform 1 0 192416 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_1770
timestamp 1694700623
transform 1 0 199584 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_1776
timestamp 1694700623
transform 1 0 200256 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_1808
timestamp 1694700623
transform 1 0 203840 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_1812
timestamp 1694700623
transform 1 0 204288 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_123_2
timestamp 1694700623
transform 1 0 1568 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_66
timestamp 1694700623
transform 1 0 8736 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_123_72
timestamp 1694700623
transform 1 0 9408 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_136
timestamp 1694700623
transform 1 0 16576 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_142
timestamp 1694700623
transform 1 0 17248 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_123_1671
timestamp 1694700623
transform 1 0 188496 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_1735
timestamp 1694700623
transform 1 0 195664 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_123_1741
timestamp 1694700623
transform 1 0 196336 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123_1805
timestamp 1694700623
transform 1 0 203504 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123_1811
timestamp 1694700623
transform 1 0 204176 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_123_1813
timestamp 1694700623
transform 1 0 204400 0 -1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_124_2
timestamp 1694700623
transform 1 0 1568 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_124_34
timestamp 1694700623
transform 1 0 5152 0 1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_124_37
timestamp 1694700623
transform 1 0 5488 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_124_101
timestamp 1694700623
transform 1 0 12656 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_124_107
timestamp 1694700623
transform 1 0 13328 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_124_139
timestamp 1694700623
transform 1 0 16912 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_143
timestamp 1694700623
transform 1 0 17360 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_124_145
timestamp 1694700623
transform 1 0 17584 0 1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_124_1671
timestamp 1694700623
transform 1 0 188496 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_124_1703
timestamp 1694700623
transform 1 0 192080 0 1 100352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_124_1706
timestamp 1694700623
transform 1 0 192416 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_124_1770
timestamp 1694700623
transform 1 0 199584 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_124_1776
timestamp 1694700623
transform 1 0 200256 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_124_1808
timestamp 1694700623
transform 1 0 203840 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124_1812
timestamp 1694700623
transform 1 0 204288 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_8
timestamp 1694700623
transform 1 0 2240 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_125_12
timestamp 1694700623
transform 1 0 2688 0 -1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_125_44
timestamp 1694700623
transform 1 0 6272 0 -1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_125_60
timestamp 1694700623
transform 1 0 8064 0 -1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_68
timestamp 1694700623
transform 1 0 8960 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_125_72
timestamp 1694700623
transform 1 0 9408 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_136
timestamp 1694700623
transform 1 0 16576 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_142
timestamp 1694700623
transform 1 0 17248 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_125_1671
timestamp 1694700623
transform 1 0 188496 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_1735
timestamp 1694700623
transform 1 0 195664 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_125_1741
timestamp 1694700623
transform 1 0 196336 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_125_1805
timestamp 1694700623
transform 1 0 203504 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_125_1811
timestamp 1694700623
transform 1 0 204176 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_125_1813
timestamp 1694700623
transform 1 0 204400 0 -1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_126_2
timestamp 1694700623
transform 1 0 1568 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_126_34
timestamp 1694700623
transform 1 0 5152 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_126_37
timestamp 1694700623
transform 1 0 5488 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_101
timestamp 1694700623
transform 1 0 12656 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_126_107
timestamp 1694700623
transform 1 0 13328 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_139
timestamp 1694700623
transform 1 0 16912 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_143
timestamp 1694700623
transform 1 0 17360 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_126_145
timestamp 1694700623
transform 1 0 17584 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_126_1671
timestamp 1694700623
transform 1 0 188496 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_126_1703
timestamp 1694700623
transform 1 0 192080 0 1 101920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_126_1706
timestamp 1694700623
transform 1 0 192416 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_126_1770
timestamp 1694700623
transform 1 0 199584 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_126_1776
timestamp 1694700623
transform 1 0 200256 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126_1808
timestamp 1694700623
transform 1 0 203840 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_127_2
timestamp 1694700623
transform 1 0 1568 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_127_66
timestamp 1694700623
transform 1 0 8736 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_127_72
timestamp 1694700623
transform 1 0 9408 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_127_136
timestamp 1694700623
transform 1 0 16576 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_127_142
timestamp 1694700623
transform 1 0 17248 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_127_1671
timestamp 1694700623
transform 1 0 188496 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_127_1735
timestamp 1694700623
transform 1 0 195664 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_127_1741
timestamp 1694700623
transform 1 0 196336 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_127_1805
timestamp 1694700623
transform 1 0 203504 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127_1811
timestamp 1694700623
transform 1 0 204176 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_127_1813
timestamp 1694700623
transform 1 0 204400 0 -1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_128_2
timestamp 1694700623
transform 1 0 1568 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_34
timestamp 1694700623
transform 1 0 5152 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_128_37
timestamp 1694700623
transform 1 0 5488 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_101
timestamp 1694700623
transform 1 0 12656 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_128_107
timestamp 1694700623
transform 1 0 13328 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_139
timestamp 1694700623
transform 1 0 16912 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_143
timestamp 1694700623
transform 1 0 17360 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_145
timestamp 1694700623
transform 1 0 17584 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_128_1671
timestamp 1694700623
transform 1 0 188496 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_128_1703
timestamp 1694700623
transform 1 0 192080 0 1 103488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_128_1706
timestamp 1694700623
transform 1 0 192416 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_1770
timestamp 1694700623
transform 1 0 199584 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_128_1776
timestamp 1694700623
transform 1 0 200256 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128_1808
timestamp 1694700623
transform 1 0 203840 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128_1812
timestamp 1694700623
transform 1 0 204288 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_129_2
timestamp 1694700623
transform 1 0 1568 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_66
timestamp 1694700623
transform 1 0 8736 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_129_72
timestamp 1694700623
transform 1 0 9408 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_136
timestamp 1694700623
transform 1 0 16576 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_142
timestamp 1694700623
transform 1 0 17248 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_129_1671
timestamp 1694700623
transform 1 0 188496 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_1735
timestamp 1694700623
transform 1 0 195664 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_129_1741
timestamp 1694700623
transform 1 0 196336 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129_1805
timestamp 1694700623
transform 1 0 203504 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129_1811
timestamp 1694700623
transform 1 0 204176 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129_1813
timestamp 1694700623
transform 1 0 204400 0 -1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_130_6
timestamp 1694700623
transform 1 0 2016 0 1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_130_22
timestamp 1694700623
transform 1 0 3808 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_30
timestamp 1694700623
transform 1 0 4704 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_34
timestamp 1694700623
transform 1 0 5152 0 1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_130_37
timestamp 1694700623
transform 1 0 5488 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_101
timestamp 1694700623
transform 1 0 12656 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_130_107
timestamp 1694700623
transform 1 0 13328 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_139
timestamp 1694700623
transform 1 0 16912 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_143
timestamp 1694700623
transform 1 0 17360 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_145
timestamp 1694700623
transform 1 0 17584 0 1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_130_1671
timestamp 1694700623
transform 1 0 188496 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130_1703
timestamp 1694700623
transform 1 0 192080 0 1 105056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_130_1706
timestamp 1694700623
transform 1 0 192416 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_1770
timestamp 1694700623
transform 1 0 199584 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_130_1776
timestamp 1694700623
transform 1 0 200256 0 1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_130_1808
timestamp 1694700623
transform 1 0 203840 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130_1812
timestamp 1694700623
transform 1 0 204288 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_131_2
timestamp 1694700623
transform 1 0 1568 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_131_66
timestamp 1694700623
transform 1 0 8736 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_131_72
timestamp 1694700623
transform 1 0 9408 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_131_136
timestamp 1694700623
transform 1 0 16576 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_131_142
timestamp 1694700623
transform 1 0 17248 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_131_1671
timestamp 1694700623
transform 1 0 188496 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_131_1735
timestamp 1694700623
transform 1 0 195664 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_131_1741
timestamp 1694700623
transform 1 0 196336 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_131_1805
timestamp 1694700623
transform 1 0 203504 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_131_1811
timestamp 1694700623
transform 1 0 204176 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_131_1813
timestamp 1694700623
transform 1 0 204400 0 -1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_132_2
timestamp 1694700623
transform 1 0 1568 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_132_34
timestamp 1694700623
transform 1 0 5152 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_132_37
timestamp 1694700623
transform 1 0 5488 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_132_101
timestamp 1694700623
transform 1 0 12656 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_132_107
timestamp 1694700623
transform 1 0 13328 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_132_139
timestamp 1694700623
transform 1 0 16912 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_143
timestamp 1694700623
transform 1 0 17360 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_132_145
timestamp 1694700623
transform 1 0 17584 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_132_1671
timestamp 1694700623
transform 1 0 188496 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_132_1703
timestamp 1694700623
transform 1 0 192080 0 1 106624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_132_1706
timestamp 1694700623
transform 1 0 192416 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_132_1770
timestamp 1694700623
transform 1 0 199584 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_132_1776
timestamp 1694700623
transform 1 0 200256 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_132_1808
timestamp 1694700623
transform 1 0 203840 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_132_1812
timestamp 1694700623
transform 1 0 204288 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_133_2
timestamp 1694700623
transform 1 0 1568 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_66
timestamp 1694700623
transform 1 0 8736 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_133_72
timestamp 1694700623
transform 1 0 9408 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_136
timestamp 1694700623
transform 1 0 16576 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_142
timestamp 1694700623
transform 1 0 17248 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_133_1671
timestamp 1694700623
transform 1 0 188496 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_1735
timestamp 1694700623
transform 1 0 195664 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_133_1741
timestamp 1694700623
transform 1 0 196336 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133_1805
timestamp 1694700623
transform 1 0 203504 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133_1811
timestamp 1694700623
transform 1 0 204176 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_133_1813
timestamp 1694700623
transform 1 0 204400 0 -1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_134_6
timestamp 1694700623
transform 1 0 2016 0 1 108192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_134_22
timestamp 1694700623
transform 1 0 3808 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_30
timestamp 1694700623
transform 1 0 4704 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_34
timestamp 1694700623
transform 1 0 5152 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_134_37
timestamp 1694700623
transform 1 0 5488 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_101
timestamp 1694700623
transform 1 0 12656 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_134_107
timestamp 1694700623
transform 1 0 13328 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_139
timestamp 1694700623
transform 1 0 16912 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_143
timestamp 1694700623
transform 1 0 17360 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_145
timestamp 1694700623
transform 1 0 17584 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_134_1671
timestamp 1694700623
transform 1 0 188496 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_134_1703
timestamp 1694700623
transform 1 0 192080 0 1 108192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_134_1706
timestamp 1694700623
transform 1 0 192416 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_1770
timestamp 1694700623
transform 1 0 199584 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_134_1776
timestamp 1694700623
transform 1 0 200256 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_134_1808
timestamp 1694700623
transform 1 0 203840 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134_1812
timestamp 1694700623
transform 1 0 204288 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_135_2
timestamp 1694700623
transform 1 0 1568 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_66
timestamp 1694700623
transform 1 0 8736 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_135_72
timestamp 1694700623
transform 1 0 9408 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_136
timestamp 1694700623
transform 1 0 16576 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_142
timestamp 1694700623
transform 1 0 17248 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_135_1671
timestamp 1694700623
transform 1 0 188496 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_1735
timestamp 1694700623
transform 1 0 195664 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_135_1741
timestamp 1694700623
transform 1 0 196336 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_135_1805
timestamp 1694700623
transform 1 0 203504 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135_1811
timestamp 1694700623
transform 1 0 204176 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135_1813
timestamp 1694700623
transform 1 0 204400 0 -1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_136_2
timestamp 1694700623
transform 1 0 1568 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_34
timestamp 1694700623
transform 1 0 5152 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_136_37
timestamp 1694700623
transform 1 0 5488 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136_101
timestamp 1694700623
transform 1 0 12656 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_136_107
timestamp 1694700623
transform 1 0 13328 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136_139
timestamp 1694700623
transform 1 0 16912 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_136_143
timestamp 1694700623
transform 1 0 17360 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_145
timestamp 1694700623
transform 1 0 17584 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_136_1671
timestamp 1694700623
transform 1 0 188496 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_136_1703
timestamp 1694700623
transform 1 0 192080 0 1 109760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_136_1706
timestamp 1694700623
transform 1 0 192416 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136_1770
timestamp 1694700623
transform 1 0 199584 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_136_1776
timestamp 1694700623
transform 1 0 200256 0 1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136_1808
timestamp 1694700623
transform 1 0 203840 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_136_1812
timestamp 1694700623
transform 1 0 204288 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_137_2
timestamp 1694700623
transform 1 0 1568 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_66
timestamp 1694700623
transform 1 0 8736 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_137_72
timestamp 1694700623
transform 1 0 9408 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_136
timestamp 1694700623
transform 1 0 16576 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_142
timestamp 1694700623
transform 1 0 17248 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_137_1671
timestamp 1694700623
transform 1 0 188496 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_1735
timestamp 1694700623
transform 1 0 195664 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_137_1741
timestamp 1694700623
transform 1 0 196336 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_137_1805
timestamp 1694700623
transform 1 0 203504 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137_1811
timestamp 1694700623
transform 1 0 204176 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_137_1813
timestamp 1694700623
transform 1 0 204400 0 -1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_2
timestamp 1694700623
transform 1 0 1568 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_138_6
timestamp 1694700623
transform 1 0 2016 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_138_22
timestamp 1694700623
transform 1 0 3808 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_30
timestamp 1694700623
transform 1 0 4704 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_34
timestamp 1694700623
transform 1 0 5152 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_138_37
timestamp 1694700623
transform 1 0 5488 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_101
timestamp 1694700623
transform 1 0 12656 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138_107
timestamp 1694700623
transform 1 0 13328 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_139
timestamp 1694700623
transform 1 0 16912 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_143
timestamp 1694700623
transform 1 0 17360 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_145
timestamp 1694700623
transform 1 0 17584 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138_1671
timestamp 1694700623
transform 1 0 188496 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_138_1703
timestamp 1694700623
transform 1 0 192080 0 1 111328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_138_1706
timestamp 1694700623
transform 1 0 192416 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_1770
timestamp 1694700623
transform 1 0 199584 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138_1776
timestamp 1694700623
transform 1 0 200256 0 1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_138_1808
timestamp 1694700623
transform 1 0 203840 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138_1812
timestamp 1694700623
transform 1 0 204288 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_139_16
timestamp 1694700623
transform 1 0 3136 0 -1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_139_48
timestamp 1694700623
transform 1 0 6720 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_64
timestamp 1694700623
transform 1 0 8512 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_68
timestamp 1694700623
transform 1 0 8960 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_139_72
timestamp 1694700623
transform 1 0 9408 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_136
timestamp 1694700623
transform 1 0 16576 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_142
timestamp 1694700623
transform 1 0 17248 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_139_1671
timestamp 1694700623
transform 1 0 188496 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_1735
timestamp 1694700623
transform 1 0 195664 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_139_1741
timestamp 1694700623
transform 1 0 196336 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_139_1805
timestamp 1694700623
transform 1 0 203504 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_139_1811
timestamp 1694700623
transform 1 0 204176 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139_1813
timestamp 1694700623
transform 1 0 204400 0 -1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_140_2
timestamp 1694700623
transform 1 0 1568 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_34
timestamp 1694700623
transform 1 0 5152 0 1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_140_37
timestamp 1694700623
transform 1 0 5488 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_101
timestamp 1694700623
transform 1 0 12656 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_140_107
timestamp 1694700623
transform 1 0 13328 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_139
timestamp 1694700623
transform 1 0 16912 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_143
timestamp 1694700623
transform 1 0 17360 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_145
timestamp 1694700623
transform 1 0 17584 0 1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_140_1671
timestamp 1694700623
transform 1 0 188496 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140_1703
timestamp 1694700623
transform 1 0 192080 0 1 112896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_140_1706
timestamp 1694700623
transform 1 0 192416 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_1770
timestamp 1694700623
transform 1 0 199584 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_140_1776
timestamp 1694700623
transform 1 0 200256 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_140_1808
timestamp 1694700623
transform 1 0 203840 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_140_1812
timestamp 1694700623
transform 1 0 204288 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_141_2
timestamp 1694700623
transform 1 0 1568 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_66
timestamp 1694700623
transform 1 0 8736 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_141_72
timestamp 1694700623
transform 1 0 9408 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_136
timestamp 1694700623
transform 1 0 16576 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_142
timestamp 1694700623
transform 1 0 17248 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_141_1671
timestamp 1694700623
transform 1 0 188496 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_1735
timestamp 1694700623
transform 1 0 195664 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_141_1741
timestamp 1694700623
transform 1 0 196336 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_141_1805
timestamp 1694700623
transform 1 0 203504 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141_1811
timestamp 1694700623
transform 1 0 204176 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_141_1813
timestamp 1694700623
transform 1 0 204400 0 -1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142_2
timestamp 1694700623
transform 1 0 1568 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142_34
timestamp 1694700623
transform 1 0 5152 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_142_37
timestamp 1694700623
transform 1 0 5488 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_101
timestamp 1694700623
transform 1 0 12656 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142_107
timestamp 1694700623
transform 1 0 13328 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_139
timestamp 1694700623
transform 1 0 16912 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142_143
timestamp 1694700623
transform 1 0 17360 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142_145
timestamp 1694700623
transform 1 0 17584 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142_1671
timestamp 1694700623
transform 1 0 188496 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142_1703
timestamp 1694700623
transform 1 0 192080 0 1 114464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_142_1706
timestamp 1694700623
transform 1 0 192416 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_1770
timestamp 1694700623
transform 1 0 199584 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142_1776
timestamp 1694700623
transform 1 0 200256 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_142_1808
timestamp 1694700623
transform 1 0 203840 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142_1812
timestamp 1694700623
transform 1 0 204288 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_143_2
timestamp 1694700623
transform 1 0 1568 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_66
timestamp 1694700623
transform 1 0 8736 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_143_72
timestamp 1694700623
transform 1 0 9408 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_136
timestamp 1694700623
transform 1 0 16576 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_142
timestamp 1694700623
transform 1 0 17248 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_143_1671
timestamp 1694700623
transform 1 0 188496 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_1735
timestamp 1694700623
transform 1 0 195664 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_143_1741
timestamp 1694700623
transform 1 0 196336 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_143_1805
timestamp 1694700623
transform 1 0 203504 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_143_1811
timestamp 1694700623
transform 1 0 204176 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_143_1813
timestamp 1694700623
transform 1 0 204400 0 -1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_144_6
timestamp 1694700623
transform 1 0 2016 0 1 116032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_144_22
timestamp 1694700623
transform 1 0 3808 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_30
timestamp 1694700623
transform 1 0 4704 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_34
timestamp 1694700623
transform 1 0 5152 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_144_37
timestamp 1694700623
transform 1 0 5488 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_101
timestamp 1694700623
transform 1 0 12656 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_144_107
timestamp 1694700623
transform 1 0 13328 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_139
timestamp 1694700623
transform 1 0 16912 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_144_143
timestamp 1694700623
transform 1 0 17360 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_145
timestamp 1694700623
transform 1 0 17584 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_144_1671
timestamp 1694700623
transform 1 0 188496 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144_1703
timestamp 1694700623
transform 1 0 192080 0 1 116032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_144_1706
timestamp 1694700623
transform 1 0 192416 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_1770
timestamp 1694700623
transform 1 0 199584 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_144_1776
timestamp 1694700623
transform 1 0 200256 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144_1808
timestamp 1694700623
transform 1 0 203840 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_144_1812
timestamp 1694700623
transform 1 0 204288 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_145_2
timestamp 1694700623
transform 1 0 1568 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_66
timestamp 1694700623
transform 1 0 8736 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_145_72
timestamp 1694700623
transform 1 0 9408 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_136
timestamp 1694700623
transform 1 0 16576 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_142
timestamp 1694700623
transform 1 0 17248 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_145_1671
timestamp 1694700623
transform 1 0 188496 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_1735
timestamp 1694700623
transform 1 0 195664 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_145_1741
timestamp 1694700623
transform 1 0 196336 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_145_1805
timestamp 1694700623
transform 1 0 203504 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145_1811
timestamp 1694700623
transform 1 0 204176 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_145_1813
timestamp 1694700623
transform 1 0 204400 0 -1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_2
timestamp 1694700623
transform 1 0 1568 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_34
timestamp 1694700623
transform 1 0 5152 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_146_37
timestamp 1694700623
transform 1 0 5488 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_101
timestamp 1694700623
transform 1 0 12656 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_107
timestamp 1694700623
transform 1 0 13328 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_139
timestamp 1694700623
transform 1 0 16912 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_143
timestamp 1694700623
transform 1 0 17360 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_145
timestamp 1694700623
transform 1 0 17584 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_1671
timestamp 1694700623
transform 1 0 188496 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_146_1703
timestamp 1694700623
transform 1 0 192080 0 1 117600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_146_1706
timestamp 1694700623
transform 1 0 192416 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_1770
timestamp 1694700623
transform 1 0 199584 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_146_1776
timestamp 1694700623
transform 1 0 200256 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_146_1808
timestamp 1694700623
transform 1 0 203840 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_146_1812
timestamp 1694700623
transform 1 0 204288 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_147_2
timestamp 1694700623
transform 1 0 1568 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_66
timestamp 1694700623
transform 1 0 8736 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_147_72
timestamp 1694700623
transform 1 0 9408 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_136
timestamp 1694700623
transform 1 0 16576 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_142
timestamp 1694700623
transform 1 0 17248 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_147_1671
timestamp 1694700623
transform 1 0 188496 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_147_1735
timestamp 1694700623
transform 1 0 195664 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_147_1741
timestamp 1694700623
transform 1 0 196336 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_1805
timestamp 1694700623
transform 1 0 203504 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147_1811
timestamp 1694700623
transform 1 0 204176 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_147_1813
timestamp 1694700623
transform 1 0 204400 0 -1 119168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_148_2
timestamp 1694700623
transform 1 0 1568 0 1 119168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_34
timestamp 1694700623
transform 1 0 5152 0 1 119168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_148_37
timestamp 1694700623
transform 1 0 5488 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_101
timestamp 1694700623
transform 1 0 12656 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_148_107
timestamp 1694700623
transform 1 0 13328 0 1 119168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_139
timestamp 1694700623
transform 1 0 16912 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_148_143
timestamp 1694700623
transform 1 0 17360 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_145
timestamp 1694700623
transform 1 0 17584 0 1 119168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_148_1671
timestamp 1694700623
transform 1 0 188496 0 1 119168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148_1703
timestamp 1694700623
transform 1 0 192080 0 1 119168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_148_1706
timestamp 1694700623
transform 1 0 192416 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_1770
timestamp 1694700623
transform 1 0 199584 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_148_1776
timestamp 1694700623
transform 1 0 200256 0 1 119168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_148_1784
timestamp 1694700623
transform 1 0 201152 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_149_6
timestamp 1694700623
transform 1 0 2016 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_149_72
timestamp 1694700623
transform 1 0 9408 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_149_136
timestamp 1694700623
transform 1 0 16576 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_149_142
timestamp 1694700623
transform 1 0 17248 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_149_1671
timestamp 1694700623
transform 1 0 188496 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_149_1735
timestamp 1694700623
transform 1 0 195664 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_149_1741
timestamp 1694700623
transform 1 0 196336 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_149_1805
timestamp 1694700623
transform 1 0 203504 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_149_1811
timestamp 1694700623
transform 1 0 204176 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_149_1813
timestamp 1694700623
transform 1 0 204400 0 -1 120736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_150_2
timestamp 1694700623
transform 1 0 1568 0 1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_150_34
timestamp 1694700623
transform 1 0 5152 0 1 120736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_150_37
timestamp 1694700623
transform 1 0 5488 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150_101
timestamp 1694700623
transform 1 0 12656 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_150_107
timestamp 1694700623
transform 1 0 13328 0 1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150_139
timestamp 1694700623
transform 1 0 16912 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150_143
timestamp 1694700623
transform 1 0 17360 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_150_145
timestamp 1694700623
transform 1 0 17584 0 1 120736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_150_1671
timestamp 1694700623
transform 1 0 188496 0 1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_150_1703
timestamp 1694700623
transform 1 0 192080 0 1 120736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_150_1706
timestamp 1694700623
transform 1 0 192416 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150_1770
timestamp 1694700623
transform 1 0 199584 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_150_1776
timestamp 1694700623
transform 1 0 200256 0 1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150_1808
timestamp 1694700623
transform 1 0 203840 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150_1812
timestamp 1694700623
transform 1 0 204288 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_151_2
timestamp 1694700623
transform 1 0 1568 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_151_66
timestamp 1694700623
transform 1 0 8736 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_151_72
timestamp 1694700623
transform 1 0 9408 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_151_136
timestamp 1694700623
transform 1 0 16576 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_151_142
timestamp 1694700623
transform 1 0 17248 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_151_1671
timestamp 1694700623
transform 1 0 188496 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_151_1735
timestamp 1694700623
transform 1 0 195664 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_151_1741
timestamp 1694700623
transform 1 0 196336 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_151_1805
timestamp 1694700623
transform 1 0 203504 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_151_1811
timestamp 1694700623
transform 1 0 204176 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_151_1813
timestamp 1694700623
transform 1 0 204400 0 -1 122304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_152_2
timestamp 1694700623
transform 1 0 1568 0 1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_152_34
timestamp 1694700623
transform 1 0 5152 0 1 122304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_152_37
timestamp 1694700623
transform 1 0 5488 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_152_101
timestamp 1694700623
transform 1 0 12656 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_152_107
timestamp 1694700623
transform 1 0 13328 0 1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_152_139
timestamp 1694700623
transform 1 0 16912 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_152_143
timestamp 1694700623
transform 1 0 17360 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_152_145
timestamp 1694700623
transform 1 0 17584 0 1 122304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_152_1671
timestamp 1694700623
transform 1 0 188496 0 1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_152_1703
timestamp 1694700623
transform 1 0 192080 0 1 122304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_152_1706
timestamp 1694700623
transform 1 0 192416 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_152_1770
timestamp 1694700623
transform 1 0 199584 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_152_1776
timestamp 1694700623
transform 1 0 200256 0 1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_152_1808
timestamp 1694700623
transform 1 0 203840 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_152_1812
timestamp 1694700623
transform 1 0 204288 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_153_2
timestamp 1694700623
transform 1 0 1568 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_153_6
timestamp 1694700623
transform 1 0 2016 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_153_72
timestamp 1694700623
transform 1 0 9408 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_153_136
timestamp 1694700623
transform 1 0 16576 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_153_142
timestamp 1694700623
transform 1 0 17248 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_153_1671
timestamp 1694700623
transform 1 0 188496 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_153_1735
timestamp 1694700623
transform 1 0 195664 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_153_1741
timestamp 1694700623
transform 1 0 196336 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_153_1805
timestamp 1694700623
transform 1 0 203504 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_153_1811
timestamp 1694700623
transform 1 0 204176 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_153_1813
timestamp 1694700623
transform 1 0 204400 0 -1 123872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_154_16
timestamp 1694700623
transform 1 0 3136 0 1 123872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_154_32
timestamp 1694700623
transform 1 0 4928 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_154_34
timestamp 1694700623
transform 1 0 5152 0 1 123872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_154_37
timestamp 1694700623
transform 1 0 5488 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_154_101
timestamp 1694700623
transform 1 0 12656 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_154_107
timestamp 1694700623
transform 1 0 13328 0 1 123872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_154_139
timestamp 1694700623
transform 1 0 16912 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_154_143
timestamp 1694700623
transform 1 0 17360 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_154_145
timestamp 1694700623
transform 1 0 17584 0 1 123872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_154_1671
timestamp 1694700623
transform 1 0 188496 0 1 123872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_154_1703
timestamp 1694700623
transform 1 0 192080 0 1 123872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_154_1706
timestamp 1694700623
transform 1 0 192416 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_154_1770
timestamp 1694700623
transform 1 0 199584 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_154_1776
timestamp 1694700623
transform 1 0 200256 0 1 123872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_154_1808
timestamp 1694700623
transform 1 0 203840 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_154_1812
timestamp 1694700623
transform 1 0 204288 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_155_2
timestamp 1694700623
transform 1 0 1568 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155_66
timestamp 1694700623
transform 1 0 8736 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_155_72
timestamp 1694700623
transform 1 0 9408 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155_136
timestamp 1694700623
transform 1 0 16576 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155_142
timestamp 1694700623
transform 1 0 17248 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_155_1671
timestamp 1694700623
transform 1 0 188496 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155_1735
timestamp 1694700623
transform 1 0 195664 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_155_1741
timestamp 1694700623
transform 1 0 196336 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_155_1805
timestamp 1694700623
transform 1 0 203504 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_155_1811
timestamp 1694700623
transform 1 0 204176 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_155_1813
timestamp 1694700623
transform 1 0 204400 0 -1 125440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_156_2
timestamp 1694700623
transform 1 0 1568 0 1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_156_34
timestamp 1694700623
transform 1 0 5152 0 1 125440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_156_37
timestamp 1694700623
transform 1 0 5488 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_156_101
timestamp 1694700623
transform 1 0 12656 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_156_107
timestamp 1694700623
transform 1 0 13328 0 1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_156_139
timestamp 1694700623
transform 1 0 16912 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_156_143
timestamp 1694700623
transform 1 0 17360 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_156_145
timestamp 1694700623
transform 1 0 17584 0 1 125440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_156_1671
timestamp 1694700623
transform 1 0 188496 0 1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_156_1703
timestamp 1694700623
transform 1 0 192080 0 1 125440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_156_1706
timestamp 1694700623
transform 1 0 192416 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_156_1770
timestamp 1694700623
transform 1 0 199584 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_156_1776
timestamp 1694700623
transform 1 0 200256 0 1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_156_1808
timestamp 1694700623
transform 1 0 203840 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_156_1812
timestamp 1694700623
transform 1 0 204288 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_157_2
timestamp 1694700623
transform 1 0 1568 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_157_66
timestamp 1694700623
transform 1 0 8736 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_157_72
timestamp 1694700623
transform 1 0 9408 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_157_136
timestamp 1694700623
transform 1 0 16576 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_157_142
timestamp 1694700623
transform 1 0 17248 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_157_1671
timestamp 1694700623
transform 1 0 188496 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_157_1735
timestamp 1694700623
transform 1 0 195664 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_157_1741
timestamp 1694700623
transform 1 0 196336 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_157_1805
timestamp 1694700623
transform 1 0 203504 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_157_1811
timestamp 1694700623
transform 1 0 204176 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_157_1813
timestamp 1694700623
transform 1 0 204400 0 -1 127008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_158_2
timestamp 1694700623
transform 1 0 1568 0 1 127008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_158_34
timestamp 1694700623
transform 1 0 5152 0 1 127008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_158_37
timestamp 1694700623
transform 1 0 5488 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158_101
timestamp 1694700623
transform 1 0 12656 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_158_107
timestamp 1694700623
transform 1 0 13328 0 1 127008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158_139
timestamp 1694700623
transform 1 0 16912 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_158_143
timestamp 1694700623
transform 1 0 17360 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_158_145
timestamp 1694700623
transform 1 0 17584 0 1 127008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_158_1671
timestamp 1694700623
transform 1 0 188496 0 1 127008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_158_1703
timestamp 1694700623
transform 1 0 192080 0 1 127008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_158_1706
timestamp 1694700623
transform 1 0 192416 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158_1770
timestamp 1694700623
transform 1 0 199584 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_158_1776
timestamp 1694700623
transform 1 0 200256 0 1 127008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_158_1808
timestamp 1694700623
transform 1 0 203840 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_158_1812
timestamp 1694700623
transform 1 0 204288 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_159_6
timestamp 1694700623
transform 1 0 2016 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_159_72
timestamp 1694700623
transform 1 0 9408 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_159_136
timestamp 1694700623
transform 1 0 16576 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_159_142
timestamp 1694700623
transform 1 0 17248 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_159_1671
timestamp 1694700623
transform 1 0 188496 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_159_1735
timestamp 1694700623
transform 1 0 195664 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_159_1741
timestamp 1694700623
transform 1 0 196336 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159_1811
timestamp 1694700623
transform 1 0 204176 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_159_1813
timestamp 1694700623
transform 1 0 204400 0 -1 128576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_160_2
timestamp 1694700623
transform 1 0 1568 0 1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_160_34
timestamp 1694700623
transform 1 0 5152 0 1 128576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_160_37
timestamp 1694700623
transform 1 0 5488 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_160_101
timestamp 1694700623
transform 1 0 12656 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_160_107
timestamp 1694700623
transform 1 0 13328 0 1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_160_139
timestamp 1694700623
transform 1 0 16912 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_160_143
timestamp 1694700623
transform 1 0 17360 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_160_145
timestamp 1694700623
transform 1 0 17584 0 1 128576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_160_1671
timestamp 1694700623
transform 1 0 188496 0 1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_160_1703
timestamp 1694700623
transform 1 0 192080 0 1 128576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_160_1706
timestamp 1694700623
transform 1 0 192416 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_160_1770
timestamp 1694700623
transform 1 0 199584 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_160_1776
timestamp 1694700623
transform 1 0 200256 0 1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_160_1808
timestamp 1694700623
transform 1 0 203840 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_160_1812
timestamp 1694700623
transform 1 0 204288 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_161_2
timestamp 1694700623
transform 1 0 1568 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_161_66
timestamp 1694700623
transform 1 0 8736 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_161_72
timestamp 1694700623
transform 1 0 9408 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_161_136
timestamp 1694700623
transform 1 0 16576 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_161_142
timestamp 1694700623
transform 1 0 17248 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_161_1671
timestamp 1694700623
transform 1 0 188496 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_161_1735
timestamp 1694700623
transform 1 0 195664 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_161_1741
timestamp 1694700623
transform 1 0 196336 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_161_1805
timestamp 1694700623
transform 1 0 203504 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_161_1811
timestamp 1694700623
transform 1 0 204176 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_161_1813
timestamp 1694700623
transform 1 0 204400 0 -1 130144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_162_2
timestamp 1694700623
transform 1 0 1568 0 1 130144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_162_34
timestamp 1694700623
transform 1 0 5152 0 1 130144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_162_37
timestamp 1694700623
transform 1 0 5488 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_162_101
timestamp 1694700623
transform 1 0 12656 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_162_107
timestamp 1694700623
transform 1 0 13328 0 1 130144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_162_139
timestamp 1694700623
transform 1 0 16912 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_162_143
timestamp 1694700623
transform 1 0 17360 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_162_145
timestamp 1694700623
transform 1 0 17584 0 1 130144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_162_1671
timestamp 1694700623
transform 1 0 188496 0 1 130144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_162_1703
timestamp 1694700623
transform 1 0 192080 0 1 130144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_162_1706
timestamp 1694700623
transform 1 0 192416 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_162_1770
timestamp 1694700623
transform 1 0 199584 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_162_1776
timestamp 1694700623
transform 1 0 200256 0 1 130144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_162_1808
timestamp 1694700623
transform 1 0 203840 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_162_1812
timestamp 1694700623
transform 1 0 204288 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_163_2
timestamp 1694700623
transform 1 0 1568 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_163_66
timestamp 1694700623
transform 1 0 8736 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_163_72
timestamp 1694700623
transform 1 0 9408 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_163_136
timestamp 1694700623
transform 1 0 16576 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_163_142
timestamp 1694700623
transform 1 0 17248 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_163_1671
timestamp 1694700623
transform 1 0 188496 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_163_1735
timestamp 1694700623
transform 1 0 195664 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_163_1741
timestamp 1694700623
transform 1 0 196336 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_163_1805
timestamp 1694700623
transform 1 0 203504 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_163_1811
timestamp 1694700623
transform 1 0 204176 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_163_1813
timestamp 1694700623
transform 1 0 204400 0 -1 131712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_164_6
timestamp 1694700623
transform 1 0 2016 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_164_22
timestamp 1694700623
transform 1 0 3808 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_164_30
timestamp 1694700623
transform 1 0 4704 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_164_34
timestamp 1694700623
transform 1 0 5152 0 1 131712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_164_37
timestamp 1694700623
transform 1 0 5488 0 1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_164_101
timestamp 1694700623
transform 1 0 12656 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_164_107
timestamp 1694700623
transform 1 0 13328 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_164_139
timestamp 1694700623
transform 1 0 16912 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_164_143
timestamp 1694700623
transform 1 0 17360 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_164_145
timestamp 1694700623
transform 1 0 17584 0 1 131712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_164_1671
timestamp 1694700623
transform 1 0 188496 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_164_1703
timestamp 1694700623
transform 1 0 192080 0 1 131712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_164_1706
timestamp 1694700623
transform 1 0 192416 0 1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_164_1770
timestamp 1694700623
transform 1 0 199584 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_164_1776
timestamp 1694700623
transform 1 0 200256 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_164_1808
timestamp 1694700623
transform 1 0 203840 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_164_1812
timestamp 1694700623
transform 1 0 204288 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_165_2
timestamp 1694700623
transform 1 0 1568 0 -1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_165_66
timestamp 1694700623
transform 1 0 8736 0 -1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_165_72
timestamp 1694700623
transform 1 0 9408 0 -1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_165_136
timestamp 1694700623
transform 1 0 16576 0 -1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_165_142
timestamp 1694700623
transform 1 0 17248 0 -1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_165_1671
timestamp 1694700623
transform 1 0 188496 0 -1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_165_1735
timestamp 1694700623
transform 1 0 195664 0 -1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_165_1741
timestamp 1694700623
transform 1 0 196336 0 -1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_165_1805
timestamp 1694700623
transform 1 0 203504 0 -1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_165_1811
timestamp 1694700623
transform 1 0 204176 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_165_1813
timestamp 1694700623
transform 1 0 204400 0 -1 133280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_166_2
timestamp 1694700623
transform 1 0 1568 0 1 133280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_166_34
timestamp 1694700623
transform 1 0 5152 0 1 133280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_166_37
timestamp 1694700623
transform 1 0 5488 0 1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_166_101
timestamp 1694700623
transform 1 0 12656 0 1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_166_107
timestamp 1694700623
transform 1 0 13328 0 1 133280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_166_139
timestamp 1694700623
transform 1 0 16912 0 1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_166_143
timestamp 1694700623
transform 1 0 17360 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_166_145
timestamp 1694700623
transform 1 0 17584 0 1 133280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_166_1671
timestamp 1694700623
transform 1 0 188496 0 1 133280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_166_1703
timestamp 1694700623
transform 1 0 192080 0 1 133280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_166_1706
timestamp 1694700623
transform 1 0 192416 0 1 133280
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_166_1770
timestamp 1694700623
transform 1 0 199584 0 1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_166_1776
timestamp 1694700623
transform 1 0 200256 0 1 133280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_166_1808
timestamp 1694700623
transform 1 0 203840 0 1 133280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_166_1812
timestamp 1694700623
transform 1 0 204288 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_167_2
timestamp 1694700623
transform 1 0 1568 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_167_6
timestamp 1694700623
transform 1 0 2016 0 -1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_167_72
timestamp 1694700623
transform 1 0 9408 0 -1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_167_136
timestamp 1694700623
transform 1 0 16576 0 -1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_167_142
timestamp 1694700623
transform 1 0 17248 0 -1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_167_1671
timestamp 1694700623
transform 1 0 188496 0 -1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_167_1735
timestamp 1694700623
transform 1 0 195664 0 -1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_167_1741
timestamp 1694700623
transform 1 0 196336 0 -1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_167_1805
timestamp 1694700623
transform 1 0 203504 0 -1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_167_1811
timestamp 1694700623
transform 1 0 204176 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_167_1813
timestamp 1694700623
transform 1 0 204400 0 -1 134848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_168_16
timestamp 1694700623
transform 1 0 3136 0 1 134848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168_32
timestamp 1694700623
transform 1 0 4928 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_168_34
timestamp 1694700623
transform 1 0 5152 0 1 134848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_168_37
timestamp 1694700623
transform 1 0 5488 0 1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_168_101
timestamp 1694700623
transform 1 0 12656 0 1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_168_107
timestamp 1694700623
transform 1 0 13328 0 1 134848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_168_139
timestamp 1694700623
transform 1 0 16912 0 1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168_143
timestamp 1694700623
transform 1 0 17360 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_168_145
timestamp 1694700623
transform 1 0 17584 0 1 134848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_168_1671
timestamp 1694700623
transform 1 0 188496 0 1 134848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_168_1703
timestamp 1694700623
transform 1 0 192080 0 1 134848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_168_1706
timestamp 1694700623
transform 1 0 192416 0 1 134848
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_168_1770
timestamp 1694700623
transform 1 0 199584 0 1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_168_1776
timestamp 1694700623
transform 1 0 200256 0 1 134848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_168_1808
timestamp 1694700623
transform 1 0 203840 0 1 134848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168_1812
timestamp 1694700623
transform 1 0 204288 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_169_2
timestamp 1694700623
transform 1 0 1568 0 -1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169_66
timestamp 1694700623
transform 1 0 8736 0 -1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_169_72
timestamp 1694700623
transform 1 0 9408 0 -1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169_136
timestamp 1694700623
transform 1 0 16576 0 -1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169_142
timestamp 1694700623
transform 1 0 17248 0 -1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_169_1671
timestamp 1694700623
transform 1 0 188496 0 -1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169_1735
timestamp 1694700623
transform 1 0 195664 0 -1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_169_1741
timestamp 1694700623
transform 1 0 196336 0 -1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169_1805
timestamp 1694700623
transform 1 0 203504 0 -1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_169_1811
timestamp 1694700623
transform 1 0 204176 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_169_1813
timestamp 1694700623
transform 1 0 204400 0 -1 136416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_170_2
timestamp 1694700623
transform 1 0 1568 0 1 136416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_170_34
timestamp 1694700623
transform 1 0 5152 0 1 136416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_170_37
timestamp 1694700623
transform 1 0 5488 0 1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_170_101
timestamp 1694700623
transform 1 0 12656 0 1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_170_107
timestamp 1694700623
transform 1 0 13328 0 1 136416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_170_139
timestamp 1694700623
transform 1 0 16912 0 1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_170_143
timestamp 1694700623
transform 1 0 17360 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_170_145
timestamp 1694700623
transform 1 0 17584 0 1 136416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_170_1671
timestamp 1694700623
transform 1 0 188496 0 1 136416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_170_1703
timestamp 1694700623
transform 1 0 192080 0 1 136416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_170_1706
timestamp 1694700623
transform 1 0 192416 0 1 136416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_170_1770
timestamp 1694700623
transform 1 0 199584 0 1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_170_1776
timestamp 1694700623
transform 1 0 200256 0 1 136416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_170_1808
timestamp 1694700623
transform 1 0 203840 0 1 136416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_170_1812
timestamp 1694700623
transform 1 0 204288 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_171_2
timestamp 1694700623
transform 1 0 1568 0 -1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171_66
timestamp 1694700623
transform 1 0 8736 0 -1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_171_72
timestamp 1694700623
transform 1 0 9408 0 -1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171_136
timestamp 1694700623
transform 1 0 16576 0 -1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171_142
timestamp 1694700623
transform 1 0 17248 0 -1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_171_1671
timestamp 1694700623
transform 1 0 188496 0 -1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171_1735
timestamp 1694700623
transform 1 0 195664 0 -1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_171_1741
timestamp 1694700623
transform 1 0 196336 0 -1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171_1805
timestamp 1694700623
transform 1 0 203504 0 -1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_171_1811
timestamp 1694700623
transform 1 0 204176 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_171_1813
timestamp 1694700623
transform 1 0 204400 0 -1 137984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172_2
timestamp 1694700623
transform 1 0 1568 0 1 137984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_172_34
timestamp 1694700623
transform 1 0 5152 0 1 137984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_172_37
timestamp 1694700623
transform 1 0 5488 0 1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_172_101
timestamp 1694700623
transform 1 0 12656 0 1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172_107
timestamp 1694700623
transform 1 0 13328 0 1 137984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_172_139
timestamp 1694700623
transform 1 0 16912 0 1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172_143
timestamp 1694700623
transform 1 0 17360 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_172_145
timestamp 1694700623
transform 1 0 17584 0 1 137984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172_1671
timestamp 1694700623
transform 1 0 188496 0 1 137984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_172_1703
timestamp 1694700623
transform 1 0 192080 0 1 137984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_172_1706
timestamp 1694700623
transform 1 0 192416 0 1 137984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_172_1770
timestamp 1694700623
transform 1 0 199584 0 1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172_1776
timestamp 1694700623
transform 1 0 200256 0 1 137984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_172_1808
timestamp 1694700623
transform 1 0 203840 0 1 137984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_172_1812
timestamp 1694700623
transform 1 0 204288 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_173_6
timestamp 1694700623
transform 1 0 2016 0 -1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_173_72
timestamp 1694700623
transform 1 0 9408 0 -1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_173_136
timestamp 1694700623
transform 1 0 16576 0 -1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_173_142
timestamp 1694700623
transform 1 0 17248 0 -1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_173_1671
timestamp 1694700623
transform 1 0 188496 0 -1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_173_1735
timestamp 1694700623
transform 1 0 195664 0 -1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_173_1741
timestamp 1694700623
transform 1 0 196336 0 -1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_173_1805
timestamp 1694700623
transform 1 0 203504 0 -1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173_1811
timestamp 1694700623
transform 1 0 204176 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_173_1813
timestamp 1694700623
transform 1 0 204400 0 -1 139552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_174_2
timestamp 1694700623
transform 1 0 1568 0 1 139552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174_34
timestamp 1694700623
transform 1 0 5152 0 1 139552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_174_37
timestamp 1694700623
transform 1 0 5488 0 1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_174_101
timestamp 1694700623
transform 1 0 12656 0 1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_174_107
timestamp 1694700623
transform 1 0 13328 0 1 139552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_174_139
timestamp 1694700623
transform 1 0 16912 0 1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_174_143
timestamp 1694700623
transform 1 0 17360 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174_145
timestamp 1694700623
transform 1 0 17584 0 1 139552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_174_1671
timestamp 1694700623
transform 1 0 188496 0 1 139552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174_1703
timestamp 1694700623
transform 1 0 192080 0 1 139552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_174_1706
timestamp 1694700623
transform 1 0 192416 0 1 139552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_174_1770
timestamp 1694700623
transform 1 0 199584 0 1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_174_1776
timestamp 1694700623
transform 1 0 200256 0 1 139552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_174_1808
timestamp 1694700623
transform 1 0 203840 0 1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_174_1812
timestamp 1694700623
transform 1 0 204288 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_175_2
timestamp 1694700623
transform 1 0 1568 0 -1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_175_66
timestamp 1694700623
transform 1 0 8736 0 -1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_175_72
timestamp 1694700623
transform 1 0 9408 0 -1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_175_136
timestamp 1694700623
transform 1 0 16576 0 -1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_175_142
timestamp 1694700623
transform 1 0 17248 0 -1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_175_1671
timestamp 1694700623
transform 1 0 188496 0 -1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_175_1735
timestamp 1694700623
transform 1 0 195664 0 -1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_175_1741
timestamp 1694700623
transform 1 0 196336 0 -1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_175_1805
timestamp 1694700623
transform 1 0 203504 0 -1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_175_1811
timestamp 1694700623
transform 1 0 204176 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_175_1813
timestamp 1694700623
transform 1 0 204400 0 -1 141120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_176_2
timestamp 1694700623
transform 1 0 1568 0 1 141120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_176_34
timestamp 1694700623
transform 1 0 5152 0 1 141120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_176_37
timestamp 1694700623
transform 1 0 5488 0 1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_176_101
timestamp 1694700623
transform 1 0 12656 0 1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_176_107
timestamp 1694700623
transform 1 0 13328 0 1 141120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_176_139
timestamp 1694700623
transform 1 0 16912 0 1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_176_143
timestamp 1694700623
transform 1 0 17360 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_176_145
timestamp 1694700623
transform 1 0 17584 0 1 141120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_176_1671
timestamp 1694700623
transform 1 0 188496 0 1 141120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_176_1703
timestamp 1694700623
transform 1 0 192080 0 1 141120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_176_1706
timestamp 1694700623
transform 1 0 192416 0 1 141120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_176_1770
timestamp 1694700623
transform 1 0 199584 0 1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_176_1776
timestamp 1694700623
transform 1 0 200256 0 1 141120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_176_1808
timestamp 1694700623
transform 1 0 203840 0 1 141120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_176_1812
timestamp 1694700623
transform 1 0 204288 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_177_2
timestamp 1694700623
transform 1 0 1568 0 -1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177_66
timestamp 1694700623
transform 1 0 8736 0 -1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_177_72
timestamp 1694700623
transform 1 0 9408 0 -1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177_136
timestamp 1694700623
transform 1 0 16576 0 -1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177_142
timestamp 1694700623
transform 1 0 17248 0 -1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_177_1671
timestamp 1694700623
transform 1 0 188496 0 -1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177_1735
timestamp 1694700623
transform 1 0 195664 0 -1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_177_1741
timestamp 1694700623
transform 1 0 196336 0 -1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177_1805
timestamp 1694700623
transform 1 0 203504 0 -1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177_1811
timestamp 1694700623
transform 1 0 204176 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177_1813
timestamp 1694700623
transform 1 0 204400 0 -1 142688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_178_6
timestamp 1694700623
transform 1 0 2016 0 1 142688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_178_22
timestamp 1694700623
transform 1 0 3808 0 1 142688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_178_30
timestamp 1694700623
transform 1 0 4704 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_178_34
timestamp 1694700623
transform 1 0 5152 0 1 142688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_178_37
timestamp 1694700623
transform 1 0 5488 0 1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_178_101
timestamp 1694700623
transform 1 0 12656 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_178_107
timestamp 1694700623
transform 1 0 13328 0 1 142688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_178_139
timestamp 1694700623
transform 1 0 16912 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_178_143
timestamp 1694700623
transform 1 0 17360 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_178_145
timestamp 1694700623
transform 1 0 17584 0 1 142688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_178_1671
timestamp 1694700623
transform 1 0 188496 0 1 142688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_178_1703
timestamp 1694700623
transform 1 0 192080 0 1 142688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_178_1706
timestamp 1694700623
transform 1 0 192416 0 1 142688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_178_1770
timestamp 1694700623
transform 1 0 199584 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_178_1776
timestamp 1694700623
transform 1 0 200256 0 1 142688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_178_1808
timestamp 1694700623
transform 1 0 203840 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_178_1812
timestamp 1694700623
transform 1 0 204288 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_179_2
timestamp 1694700623
transform 1 0 1568 0 -1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_179_66
timestamp 1694700623
transform 1 0 8736 0 -1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_179_72
timestamp 1694700623
transform 1 0 9408 0 -1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_179_136
timestamp 1694700623
transform 1 0 16576 0 -1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_179_142
timestamp 1694700623
transform 1 0 17248 0 -1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_179_1671
timestamp 1694700623
transform 1 0 188496 0 -1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_179_1735
timestamp 1694700623
transform 1 0 195664 0 -1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_179_1741
timestamp 1694700623
transform 1 0 196336 0 -1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_179_1805
timestamp 1694700623
transform 1 0 203504 0 -1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_179_1811
timestamp 1694700623
transform 1 0 204176 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_179_1813
timestamp 1694700623
transform 1 0 204400 0 -1 144256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_180_2
timestamp 1694700623
transform 1 0 1568 0 1 144256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_180_34
timestamp 1694700623
transform 1 0 5152 0 1 144256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_180_37
timestamp 1694700623
transform 1 0 5488 0 1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_180_101
timestamp 1694700623
transform 1 0 12656 0 1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_180_107
timestamp 1694700623
transform 1 0 13328 0 1 144256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_180_139
timestamp 1694700623
transform 1 0 16912 0 1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_180_143
timestamp 1694700623
transform 1 0 17360 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_180_145
timestamp 1694700623
transform 1 0 17584 0 1 144256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_180_1671
timestamp 1694700623
transform 1 0 188496 0 1 144256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_180_1703
timestamp 1694700623
transform 1 0 192080 0 1 144256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_180_1706
timestamp 1694700623
transform 1 0 192416 0 1 144256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_180_1770
timestamp 1694700623
transform 1 0 199584 0 1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_180_1776
timestamp 1694700623
transform 1 0 200256 0 1 144256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_180_1808
timestamp 1694700623
transform 1 0 203840 0 1 144256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_180_1812
timestamp 1694700623
transform 1 0 204288 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_2
timestamp 1694700623
transform 1 0 1568 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_36
timestamp 1694700623
transform 1 0 5376 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_70
timestamp 1694700623
transform 1 0 9184 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_104
timestamp 1694700623
transform 1 0 12992 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_138
timestamp 1694700623
transform 1 0 16800 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_172
timestamp 1694700623
transform 1 0 20608 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_206
timestamp 1694700623
transform 1 0 24416 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_240
timestamp 1694700623
transform 1 0 28224 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_274
timestamp 1694700623
transform 1 0 32032 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_308
timestamp 1694700623
transform 1 0 35840 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_342
timestamp 1694700623
transform 1 0 39648 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_376
timestamp 1694700623
transform 1 0 43456 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_410
timestamp 1694700623
transform 1 0 47264 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_444
timestamp 1694700623
transform 1 0 51072 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_478
timestamp 1694700623
transform 1 0 54880 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_512
timestamp 1694700623
transform 1 0 58688 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_546
timestamp 1694700623
transform 1 0 62496 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_580
timestamp 1694700623
transform 1 0 66304 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_614
timestamp 1694700623
transform 1 0 70112 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_648
timestamp 1694700623
transform 1 0 73920 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_682
timestamp 1694700623
transform 1 0 77728 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_716
timestamp 1694700623
transform 1 0 81536 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_750
timestamp 1694700623
transform 1 0 85344 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_784
timestamp 1694700623
transform 1 0 89152 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_818
timestamp 1694700623
transform 1 0 92960 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_852
timestamp 1694700623
transform 1 0 96768 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_886
timestamp 1694700623
transform 1 0 100576 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_920
timestamp 1694700623
transform 1 0 104384 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_954
timestamp 1694700623
transform 1 0 108192 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_988
timestamp 1694700623
transform 1 0 112000 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1022
timestamp 1694700623
transform 1 0 115808 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1056
timestamp 1694700623
transform 1 0 119616 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1090
timestamp 1694700623
transform 1 0 123424 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1124
timestamp 1694700623
transform 1 0 127232 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1158
timestamp 1694700623
transform 1 0 131040 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1192
timestamp 1694700623
transform 1 0 134848 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1226
timestamp 1694700623
transform 1 0 138656 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1260
timestamp 1694700623
transform 1 0 142464 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1294
timestamp 1694700623
transform 1 0 146272 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1328
timestamp 1694700623
transform 1 0 150080 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1362
timestamp 1694700623
transform 1 0 153888 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1396
timestamp 1694700623
transform 1 0 157696 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1430
timestamp 1694700623
transform 1 0 161504 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1464
timestamp 1694700623
transform 1 0 165312 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1498
timestamp 1694700623
transform 1 0 169120 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1532
timestamp 1694700623
transform 1 0 172928 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1566
timestamp 1694700623
transform 1 0 176736 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1600
timestamp 1694700623
transform 1 0 180544 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1634
timestamp 1694700623
transform 1 0 184352 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1668
timestamp 1694700623
transform 1 0 188160 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1702
timestamp 1694700623
transform 1 0 191968 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1736
timestamp 1694700623
transform 1 0 195776 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_181_1770
timestamp 1694700623
transform 1 0 199584 0 -1 145824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_181_1804
timestamp 1694700623
transform 1 0 203392 0 -1 145824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_181_1812
timestamp 1694700623
transform 1 0 204288 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_182_2
timestamp 1694700623
transform 1 0 1568 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_182_6
timestamp 1694700623
transform 1 0 2016 0 1 145824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182_22
timestamp 1694700623
transform 1 0 3808 0 1 145824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_30
timestamp 1694700623
transform 1 0 4704 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_182_34
timestamp 1694700623
transform 1 0 5152 0 1 145824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_37
timestamp 1694700623
transform 1 0 5488 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_101
timestamp 1694700623
transform 1 0 12656 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_107
timestamp 1694700623
transform 1 0 13328 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_171
timestamp 1694700623
transform 1 0 20496 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_177
timestamp 1694700623
transform 1 0 21168 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_241
timestamp 1694700623
transform 1 0 28336 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_247
timestamp 1694700623
transform 1 0 29008 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_311
timestamp 1694700623
transform 1 0 36176 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_317
timestamp 1694700623
transform 1 0 36848 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_381
timestamp 1694700623
transform 1 0 44016 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_387
timestamp 1694700623
transform 1 0 44688 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_451
timestamp 1694700623
transform 1 0 51856 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_457
timestamp 1694700623
transform 1 0 52528 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_521
timestamp 1694700623
transform 1 0 59696 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_527
timestamp 1694700623
transform 1 0 60368 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_591
timestamp 1694700623
transform 1 0 67536 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_597
timestamp 1694700623
transform 1 0 68208 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_661
timestamp 1694700623
transform 1 0 75376 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_667
timestamp 1694700623
transform 1 0 76048 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_731
timestamp 1694700623
transform 1 0 83216 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_737
timestamp 1694700623
transform 1 0 83888 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_801
timestamp 1694700623
transform 1 0 91056 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_807
timestamp 1694700623
transform 1 0 91728 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_871
timestamp 1694700623
transform 1 0 98896 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_877
timestamp 1694700623
transform 1 0 99568 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_941
timestamp 1694700623
transform 1 0 106736 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_947
timestamp 1694700623
transform 1 0 107408 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1011
timestamp 1694700623
transform 1 0 114576 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1017
timestamp 1694700623
transform 1 0 115248 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1081
timestamp 1694700623
transform 1 0 122416 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1087
timestamp 1694700623
transform 1 0 123088 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1151
timestamp 1694700623
transform 1 0 130256 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1157
timestamp 1694700623
transform 1 0 130928 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1221
timestamp 1694700623
transform 1 0 138096 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1227
timestamp 1694700623
transform 1 0 138768 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1291
timestamp 1694700623
transform 1 0 145936 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1297
timestamp 1694700623
transform 1 0 146608 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1361
timestamp 1694700623
transform 1 0 153776 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1367
timestamp 1694700623
transform 1 0 154448 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1431
timestamp 1694700623
transform 1 0 161616 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1437
timestamp 1694700623
transform 1 0 162288 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1501
timestamp 1694700623
transform 1 0 169456 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1507
timestamp 1694700623
transform 1 0 170128 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1571
timestamp 1694700623
transform 1 0 177296 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1577
timestamp 1694700623
transform 1 0 177968 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1641
timestamp 1694700623
transform 1 0 185136 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1647
timestamp 1694700623
transform 1 0 185808 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_182_1711
timestamp 1694700623
transform 1 0 192976 0 1 145824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_182_1717
timestamp 1694700623
transform 1 0 193648 0 1 145824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_182_1781
timestamp 1694700623
transform 1 0 200816 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_182_1787
timestamp 1694700623
transform 1 0 201488 0 1 145824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_183_16
timestamp 1694700623
transform 1 0 3136 0 -1 147392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_183_48
timestamp 1694700623
transform 1 0 6720 0 -1 147392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_64
timestamp 1694700623
transform 1 0 8512 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_183_68
timestamp 1694700623
transform 1 0 8960 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_72
timestamp 1694700623
transform 1 0 9408 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_136
timestamp 1694700623
transform 1 0 16576 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_142
timestamp 1694700623
transform 1 0 17248 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_206
timestamp 1694700623
transform 1 0 24416 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_212
timestamp 1694700623
transform 1 0 25088 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_276
timestamp 1694700623
transform 1 0 32256 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_282
timestamp 1694700623
transform 1 0 32928 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_346
timestamp 1694700623
transform 1 0 40096 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_352
timestamp 1694700623
transform 1 0 40768 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_416
timestamp 1694700623
transform 1 0 47936 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_422
timestamp 1694700623
transform 1 0 48608 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_486
timestamp 1694700623
transform 1 0 55776 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_492
timestamp 1694700623
transform 1 0 56448 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_556
timestamp 1694700623
transform 1 0 63616 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_562
timestamp 1694700623
transform 1 0 64288 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_626
timestamp 1694700623
transform 1 0 71456 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_632
timestamp 1694700623
transform 1 0 72128 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_696
timestamp 1694700623
transform 1 0 79296 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_702
timestamp 1694700623
transform 1 0 79968 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_766
timestamp 1694700623
transform 1 0 87136 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_772
timestamp 1694700623
transform 1 0 87808 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_836
timestamp 1694700623
transform 1 0 94976 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_842
timestamp 1694700623
transform 1 0 95648 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_906
timestamp 1694700623
transform 1 0 102816 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_912
timestamp 1694700623
transform 1 0 103488 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_976
timestamp 1694700623
transform 1 0 110656 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_982
timestamp 1694700623
transform 1 0 111328 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1046
timestamp 1694700623
transform 1 0 118496 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1052
timestamp 1694700623
transform 1 0 119168 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1116
timestamp 1694700623
transform 1 0 126336 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1122
timestamp 1694700623
transform 1 0 127008 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1186
timestamp 1694700623
transform 1 0 134176 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1192
timestamp 1694700623
transform 1 0 134848 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1256
timestamp 1694700623
transform 1 0 142016 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1262
timestamp 1694700623
transform 1 0 142688 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1326
timestamp 1694700623
transform 1 0 149856 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1332
timestamp 1694700623
transform 1 0 150528 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1396
timestamp 1694700623
transform 1 0 157696 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1402
timestamp 1694700623
transform 1 0 158368 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1466
timestamp 1694700623
transform 1 0 165536 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1472
timestamp 1694700623
transform 1 0 166208 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1536
timestamp 1694700623
transform 1 0 173376 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1542
timestamp 1694700623
transform 1 0 174048 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1606
timestamp 1694700623
transform 1 0 181216 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1612
timestamp 1694700623
transform 1 0 181888 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1676
timestamp 1694700623
transform 1 0 189056 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_183_1682
timestamp 1694700623
transform 1 0 189728 0 -1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1746
timestamp 1694700623
transform 1 0 196896 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_183_1752
timestamp 1694700623
transform 1 0 197568 0 -1 147392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_183_1784
timestamp 1694700623
transform 1 0 201152 0 -1 147392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_183_1800
timestamp 1694700623
transform 1 0 202944 0 -1 147392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_183_1808
timestamp 1694700623
transform 1 0 203840 0 -1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_183_1812
timestamp 1694700623
transform 1 0 204288 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_184_2
timestamp 1694700623
transform 1 0 1568 0 1 147392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_184_34
timestamp 1694700623
transform 1 0 5152 0 1 147392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_37
timestamp 1694700623
transform 1 0 5488 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_101
timestamp 1694700623
transform 1 0 12656 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_107
timestamp 1694700623
transform 1 0 13328 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_171
timestamp 1694700623
transform 1 0 20496 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_177
timestamp 1694700623
transform 1 0 21168 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_241
timestamp 1694700623
transform 1 0 28336 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_247
timestamp 1694700623
transform 1 0 29008 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_311
timestamp 1694700623
transform 1 0 36176 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_317
timestamp 1694700623
transform 1 0 36848 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_381
timestamp 1694700623
transform 1 0 44016 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_387
timestamp 1694700623
transform 1 0 44688 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_451
timestamp 1694700623
transform 1 0 51856 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_457
timestamp 1694700623
transform 1 0 52528 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_521
timestamp 1694700623
transform 1 0 59696 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_527
timestamp 1694700623
transform 1 0 60368 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_591
timestamp 1694700623
transform 1 0 67536 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_597
timestamp 1694700623
transform 1 0 68208 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_661
timestamp 1694700623
transform 1 0 75376 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_667
timestamp 1694700623
transform 1 0 76048 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_731
timestamp 1694700623
transform 1 0 83216 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_737
timestamp 1694700623
transform 1 0 83888 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_801
timestamp 1694700623
transform 1 0 91056 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_807
timestamp 1694700623
transform 1 0 91728 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_871
timestamp 1694700623
transform 1 0 98896 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_877
timestamp 1694700623
transform 1 0 99568 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_941
timestamp 1694700623
transform 1 0 106736 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_947
timestamp 1694700623
transform 1 0 107408 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1011
timestamp 1694700623
transform 1 0 114576 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1017
timestamp 1694700623
transform 1 0 115248 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1081
timestamp 1694700623
transform 1 0 122416 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1087
timestamp 1694700623
transform 1 0 123088 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1151
timestamp 1694700623
transform 1 0 130256 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1157
timestamp 1694700623
transform 1 0 130928 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1221
timestamp 1694700623
transform 1 0 138096 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1227
timestamp 1694700623
transform 1 0 138768 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1291
timestamp 1694700623
transform 1 0 145936 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1297
timestamp 1694700623
transform 1 0 146608 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1361
timestamp 1694700623
transform 1 0 153776 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1367
timestamp 1694700623
transform 1 0 154448 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1431
timestamp 1694700623
transform 1 0 161616 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1437
timestamp 1694700623
transform 1 0 162288 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1501
timestamp 1694700623
transform 1 0 169456 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1507
timestamp 1694700623
transform 1 0 170128 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1571
timestamp 1694700623
transform 1 0 177296 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1577
timestamp 1694700623
transform 1 0 177968 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1641
timestamp 1694700623
transform 1 0 185136 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1647
timestamp 1694700623
transform 1 0 185808 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1711
timestamp 1694700623
transform 1 0 192976 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_184_1717
timestamp 1694700623
transform 1 0 193648 0 1 147392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_184_1781
timestamp 1694700623
transform 1 0 200816 0 1 147392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_184_1787
timestamp 1694700623
transform 1 0 201488 0 1 147392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_184_1803
timestamp 1694700623
transform 1 0 203280 0 1 147392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_184_1811
timestamp 1694700623
transform 1 0 204176 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_184_1813
timestamp 1694700623
transform 1 0 204400 0 1 147392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_2
timestamp 1694700623
transform 1 0 1568 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_66
timestamp 1694700623
transform 1 0 8736 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_72
timestamp 1694700623
transform 1 0 9408 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_136
timestamp 1694700623
transform 1 0 16576 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_142
timestamp 1694700623
transform 1 0 17248 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_206
timestamp 1694700623
transform 1 0 24416 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_212
timestamp 1694700623
transform 1 0 25088 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_276
timestamp 1694700623
transform 1 0 32256 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_282
timestamp 1694700623
transform 1 0 32928 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_346
timestamp 1694700623
transform 1 0 40096 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_352
timestamp 1694700623
transform 1 0 40768 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_416
timestamp 1694700623
transform 1 0 47936 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_422
timestamp 1694700623
transform 1 0 48608 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_486
timestamp 1694700623
transform 1 0 55776 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_492
timestamp 1694700623
transform 1 0 56448 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_556
timestamp 1694700623
transform 1 0 63616 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_562
timestamp 1694700623
transform 1 0 64288 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_626
timestamp 1694700623
transform 1 0 71456 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_632
timestamp 1694700623
transform 1 0 72128 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_696
timestamp 1694700623
transform 1 0 79296 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_702
timestamp 1694700623
transform 1 0 79968 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_766
timestamp 1694700623
transform 1 0 87136 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_772
timestamp 1694700623
transform 1 0 87808 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_836
timestamp 1694700623
transform 1 0 94976 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_842
timestamp 1694700623
transform 1 0 95648 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_906
timestamp 1694700623
transform 1 0 102816 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_912
timestamp 1694700623
transform 1 0 103488 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_976
timestamp 1694700623
transform 1 0 110656 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_982
timestamp 1694700623
transform 1 0 111328 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1046
timestamp 1694700623
transform 1 0 118496 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1052
timestamp 1694700623
transform 1 0 119168 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1116
timestamp 1694700623
transform 1 0 126336 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1122
timestamp 1694700623
transform 1 0 127008 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1186
timestamp 1694700623
transform 1 0 134176 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1192
timestamp 1694700623
transform 1 0 134848 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1256
timestamp 1694700623
transform 1 0 142016 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1262
timestamp 1694700623
transform 1 0 142688 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1326
timestamp 1694700623
transform 1 0 149856 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1332
timestamp 1694700623
transform 1 0 150528 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1396
timestamp 1694700623
transform 1 0 157696 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1402
timestamp 1694700623
transform 1 0 158368 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1466
timestamp 1694700623
transform 1 0 165536 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1472
timestamp 1694700623
transform 1 0 166208 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1536
timestamp 1694700623
transform 1 0 173376 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1542
timestamp 1694700623
transform 1 0 174048 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1606
timestamp 1694700623
transform 1 0 181216 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1612
timestamp 1694700623
transform 1 0 181888 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1676
timestamp 1694700623
transform 1 0 189056 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_185_1682
timestamp 1694700623
transform 1 0 189728 0 -1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1746
timestamp 1694700623
transform 1 0 196896 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_185_1752
timestamp 1694700623
transform 1 0 197568 0 -1 148960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_185_1784
timestamp 1694700623
transform 1 0 201152 0 -1 148960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_185_1800
timestamp 1694700623
transform 1 0 202944 0 -1 148960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_185_1808
timestamp 1694700623
transform 1 0 203840 0 -1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185_1812
timestamp 1694700623
transform 1 0 204288 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_186_2
timestamp 1694700623
transform 1 0 1568 0 1 148960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_186_34
timestamp 1694700623
transform 1 0 5152 0 1 148960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_37
timestamp 1694700623
transform 1 0 5488 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_101
timestamp 1694700623
transform 1 0 12656 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_107
timestamp 1694700623
transform 1 0 13328 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_171
timestamp 1694700623
transform 1 0 20496 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_177
timestamp 1694700623
transform 1 0 21168 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_241
timestamp 1694700623
transform 1 0 28336 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_247
timestamp 1694700623
transform 1 0 29008 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_311
timestamp 1694700623
transform 1 0 36176 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_317
timestamp 1694700623
transform 1 0 36848 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_381
timestamp 1694700623
transform 1 0 44016 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_387
timestamp 1694700623
transform 1 0 44688 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_451
timestamp 1694700623
transform 1 0 51856 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_457
timestamp 1694700623
transform 1 0 52528 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_521
timestamp 1694700623
transform 1 0 59696 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_527
timestamp 1694700623
transform 1 0 60368 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_591
timestamp 1694700623
transform 1 0 67536 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_597
timestamp 1694700623
transform 1 0 68208 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_661
timestamp 1694700623
transform 1 0 75376 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_667
timestamp 1694700623
transform 1 0 76048 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_731
timestamp 1694700623
transform 1 0 83216 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_737
timestamp 1694700623
transform 1 0 83888 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_801
timestamp 1694700623
transform 1 0 91056 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_807
timestamp 1694700623
transform 1 0 91728 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_871
timestamp 1694700623
transform 1 0 98896 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_877
timestamp 1694700623
transform 1 0 99568 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_941
timestamp 1694700623
transform 1 0 106736 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_947
timestamp 1694700623
transform 1 0 107408 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1011
timestamp 1694700623
transform 1 0 114576 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1017
timestamp 1694700623
transform 1 0 115248 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1081
timestamp 1694700623
transform 1 0 122416 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1087
timestamp 1694700623
transform 1 0 123088 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1151
timestamp 1694700623
transform 1 0 130256 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1157
timestamp 1694700623
transform 1 0 130928 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1221
timestamp 1694700623
transform 1 0 138096 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1227
timestamp 1694700623
transform 1 0 138768 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1291
timestamp 1694700623
transform 1 0 145936 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1297
timestamp 1694700623
transform 1 0 146608 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1361
timestamp 1694700623
transform 1 0 153776 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1367
timestamp 1694700623
transform 1 0 154448 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1431
timestamp 1694700623
transform 1 0 161616 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1437
timestamp 1694700623
transform 1 0 162288 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1501
timestamp 1694700623
transform 1 0 169456 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1507
timestamp 1694700623
transform 1 0 170128 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1571
timestamp 1694700623
transform 1 0 177296 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1577
timestamp 1694700623
transform 1 0 177968 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1641
timestamp 1694700623
transform 1 0 185136 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1647
timestamp 1694700623
transform 1 0 185808 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1711
timestamp 1694700623
transform 1 0 192976 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_186_1717
timestamp 1694700623
transform 1 0 193648 0 1 148960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_186_1781
timestamp 1694700623
transform 1 0 200816 0 1 148960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_186_1787
timestamp 1694700623
transform 1 0 201488 0 1 148960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_186_1803
timestamp 1694700623
transform 1 0 203280 0 1 148960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_186_1811
timestamp 1694700623
transform 1 0 204176 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_186_1813
timestamp 1694700623
transform 1 0 204400 0 1 148960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_2
timestamp 1694700623
transform 1 0 1568 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_66
timestamp 1694700623
transform 1 0 8736 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_72
timestamp 1694700623
transform 1 0 9408 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_136
timestamp 1694700623
transform 1 0 16576 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_142
timestamp 1694700623
transform 1 0 17248 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_206
timestamp 1694700623
transform 1 0 24416 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_212
timestamp 1694700623
transform 1 0 25088 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_276
timestamp 1694700623
transform 1 0 32256 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_282
timestamp 1694700623
transform 1 0 32928 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_346
timestamp 1694700623
transform 1 0 40096 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_352
timestamp 1694700623
transform 1 0 40768 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_416
timestamp 1694700623
transform 1 0 47936 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_422
timestamp 1694700623
transform 1 0 48608 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_486
timestamp 1694700623
transform 1 0 55776 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_492
timestamp 1694700623
transform 1 0 56448 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_556
timestamp 1694700623
transform 1 0 63616 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_562
timestamp 1694700623
transform 1 0 64288 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_626
timestamp 1694700623
transform 1 0 71456 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_632
timestamp 1694700623
transform 1 0 72128 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_696
timestamp 1694700623
transform 1 0 79296 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_702
timestamp 1694700623
transform 1 0 79968 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_766
timestamp 1694700623
transform 1 0 87136 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_772
timestamp 1694700623
transform 1 0 87808 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_836
timestamp 1694700623
transform 1 0 94976 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_842
timestamp 1694700623
transform 1 0 95648 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_906
timestamp 1694700623
transform 1 0 102816 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_912
timestamp 1694700623
transform 1 0 103488 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_976
timestamp 1694700623
transform 1 0 110656 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_982
timestamp 1694700623
transform 1 0 111328 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1046
timestamp 1694700623
transform 1 0 118496 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1052
timestamp 1694700623
transform 1 0 119168 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1116
timestamp 1694700623
transform 1 0 126336 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1122
timestamp 1694700623
transform 1 0 127008 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1186
timestamp 1694700623
transform 1 0 134176 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1192
timestamp 1694700623
transform 1 0 134848 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1256
timestamp 1694700623
transform 1 0 142016 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1262
timestamp 1694700623
transform 1 0 142688 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1326
timestamp 1694700623
transform 1 0 149856 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1332
timestamp 1694700623
transform 1 0 150528 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1396
timestamp 1694700623
transform 1 0 157696 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1402
timestamp 1694700623
transform 1 0 158368 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1466
timestamp 1694700623
transform 1 0 165536 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1472
timestamp 1694700623
transform 1 0 166208 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1536
timestamp 1694700623
transform 1 0 173376 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1542
timestamp 1694700623
transform 1 0 174048 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1606
timestamp 1694700623
transform 1 0 181216 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1612
timestamp 1694700623
transform 1 0 181888 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1676
timestamp 1694700623
transform 1 0 189056 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_187_1682
timestamp 1694700623
transform 1 0 189728 0 -1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1746
timestamp 1694700623
transform 1 0 196896 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_187_1752
timestamp 1694700623
transform 1 0 197568 0 -1 150528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_187_1784
timestamp 1694700623
transform 1 0 201152 0 -1 150528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_187_1800
timestamp 1694700623
transform 1 0 202944 0 -1 150528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187_1808
timestamp 1694700623
transform 1 0 203840 0 -1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_187_1812
timestamp 1694700623
transform 1 0 204288 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_188_6
timestamp 1694700623
transform 1 0 2016 0 1 150528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_188_22
timestamp 1694700623
transform 1 0 3808 0 1 150528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_30
timestamp 1694700623
transform 1 0 4704 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_188_34
timestamp 1694700623
transform 1 0 5152 0 1 150528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_37
timestamp 1694700623
transform 1 0 5488 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_101
timestamp 1694700623
transform 1 0 12656 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_107
timestamp 1694700623
transform 1 0 13328 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_171
timestamp 1694700623
transform 1 0 20496 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_177
timestamp 1694700623
transform 1 0 21168 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_241
timestamp 1694700623
transform 1 0 28336 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_247
timestamp 1694700623
transform 1 0 29008 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_311
timestamp 1694700623
transform 1 0 36176 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_317
timestamp 1694700623
transform 1 0 36848 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_381
timestamp 1694700623
transform 1 0 44016 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_387
timestamp 1694700623
transform 1 0 44688 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_451
timestamp 1694700623
transform 1 0 51856 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_457
timestamp 1694700623
transform 1 0 52528 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_521
timestamp 1694700623
transform 1 0 59696 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_527
timestamp 1694700623
transform 1 0 60368 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_591
timestamp 1694700623
transform 1 0 67536 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_597
timestamp 1694700623
transform 1 0 68208 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_661
timestamp 1694700623
transform 1 0 75376 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_667
timestamp 1694700623
transform 1 0 76048 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_731
timestamp 1694700623
transform 1 0 83216 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_737
timestamp 1694700623
transform 1 0 83888 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_801
timestamp 1694700623
transform 1 0 91056 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_807
timestamp 1694700623
transform 1 0 91728 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_871
timestamp 1694700623
transform 1 0 98896 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_877
timestamp 1694700623
transform 1 0 99568 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_941
timestamp 1694700623
transform 1 0 106736 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_947
timestamp 1694700623
transform 1 0 107408 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1011
timestamp 1694700623
transform 1 0 114576 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1017
timestamp 1694700623
transform 1 0 115248 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1081
timestamp 1694700623
transform 1 0 122416 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1087
timestamp 1694700623
transform 1 0 123088 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1151
timestamp 1694700623
transform 1 0 130256 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1157
timestamp 1694700623
transform 1 0 130928 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1221
timestamp 1694700623
transform 1 0 138096 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1227
timestamp 1694700623
transform 1 0 138768 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1291
timestamp 1694700623
transform 1 0 145936 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1297
timestamp 1694700623
transform 1 0 146608 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1361
timestamp 1694700623
transform 1 0 153776 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1367
timestamp 1694700623
transform 1 0 154448 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1431
timestamp 1694700623
transform 1 0 161616 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1437
timestamp 1694700623
transform 1 0 162288 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1501
timestamp 1694700623
transform 1 0 169456 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1507
timestamp 1694700623
transform 1 0 170128 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1571
timestamp 1694700623
transform 1 0 177296 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1577
timestamp 1694700623
transform 1 0 177968 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1641
timestamp 1694700623
transform 1 0 185136 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1647
timestamp 1694700623
transform 1 0 185808 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1711
timestamp 1694700623
transform 1 0 192976 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_188_1717
timestamp 1694700623
transform 1 0 193648 0 1 150528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188_1781
timestamp 1694700623
transform 1 0 200816 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_188_1787
timestamp 1694700623
transform 1 0 201488 0 1 150528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_188_1803
timestamp 1694700623
transform 1 0 203280 0 1 150528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_188_1811
timestamp 1694700623
transform 1 0 204176 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_188_1813
timestamp 1694700623
transform 1 0 204400 0 1 150528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_2
timestamp 1694700623
transform 1 0 1568 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_66
timestamp 1694700623
transform 1 0 8736 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_72
timestamp 1694700623
transform 1 0 9408 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_136
timestamp 1694700623
transform 1 0 16576 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_142
timestamp 1694700623
transform 1 0 17248 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_206
timestamp 1694700623
transform 1 0 24416 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_212
timestamp 1694700623
transform 1 0 25088 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_276
timestamp 1694700623
transform 1 0 32256 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_282
timestamp 1694700623
transform 1 0 32928 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_346
timestamp 1694700623
transform 1 0 40096 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_352
timestamp 1694700623
transform 1 0 40768 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_416
timestamp 1694700623
transform 1 0 47936 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_422
timestamp 1694700623
transform 1 0 48608 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_486
timestamp 1694700623
transform 1 0 55776 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_492
timestamp 1694700623
transform 1 0 56448 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_556
timestamp 1694700623
transform 1 0 63616 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_562
timestamp 1694700623
transform 1 0 64288 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_626
timestamp 1694700623
transform 1 0 71456 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_632
timestamp 1694700623
transform 1 0 72128 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_696
timestamp 1694700623
transform 1 0 79296 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_702
timestamp 1694700623
transform 1 0 79968 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_766
timestamp 1694700623
transform 1 0 87136 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_772
timestamp 1694700623
transform 1 0 87808 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_836
timestamp 1694700623
transform 1 0 94976 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_842
timestamp 1694700623
transform 1 0 95648 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_906
timestamp 1694700623
transform 1 0 102816 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_912
timestamp 1694700623
transform 1 0 103488 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_976
timestamp 1694700623
transform 1 0 110656 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_982
timestamp 1694700623
transform 1 0 111328 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1046
timestamp 1694700623
transform 1 0 118496 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1052
timestamp 1694700623
transform 1 0 119168 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1116
timestamp 1694700623
transform 1 0 126336 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1122
timestamp 1694700623
transform 1 0 127008 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1186
timestamp 1694700623
transform 1 0 134176 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1192
timestamp 1694700623
transform 1 0 134848 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1256
timestamp 1694700623
transform 1 0 142016 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1262
timestamp 1694700623
transform 1 0 142688 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1326
timestamp 1694700623
transform 1 0 149856 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1332
timestamp 1694700623
transform 1 0 150528 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1396
timestamp 1694700623
transform 1 0 157696 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1402
timestamp 1694700623
transform 1 0 158368 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1466
timestamp 1694700623
transform 1 0 165536 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1472
timestamp 1694700623
transform 1 0 166208 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1536
timestamp 1694700623
transform 1 0 173376 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1542
timestamp 1694700623
transform 1 0 174048 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1606
timestamp 1694700623
transform 1 0 181216 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1612
timestamp 1694700623
transform 1 0 181888 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1676
timestamp 1694700623
transform 1 0 189056 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_189_1682
timestamp 1694700623
transform 1 0 189728 0 -1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1746
timestamp 1694700623
transform 1 0 196896 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_189_1752
timestamp 1694700623
transform 1 0 197568 0 -1 152096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_189_1784
timestamp 1694700623
transform 1 0 201152 0 -1 152096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_189_1800
timestamp 1694700623
transform 1 0 202944 0 -1 152096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_189_1808
timestamp 1694700623
transform 1 0 203840 0 -1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_189_1812
timestamp 1694700623
transform 1 0 204288 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_190_2
timestamp 1694700623
transform 1 0 1568 0 1 152096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_190_34
timestamp 1694700623
transform 1 0 5152 0 1 152096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_37
timestamp 1694700623
transform 1 0 5488 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_101
timestamp 1694700623
transform 1 0 12656 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_107
timestamp 1694700623
transform 1 0 13328 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_171
timestamp 1694700623
transform 1 0 20496 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_177
timestamp 1694700623
transform 1 0 21168 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_241
timestamp 1694700623
transform 1 0 28336 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_247
timestamp 1694700623
transform 1 0 29008 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_311
timestamp 1694700623
transform 1 0 36176 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_317
timestamp 1694700623
transform 1 0 36848 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_381
timestamp 1694700623
transform 1 0 44016 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_387
timestamp 1694700623
transform 1 0 44688 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_451
timestamp 1694700623
transform 1 0 51856 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_457
timestamp 1694700623
transform 1 0 52528 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_521
timestamp 1694700623
transform 1 0 59696 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_527
timestamp 1694700623
transform 1 0 60368 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_591
timestamp 1694700623
transform 1 0 67536 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_597
timestamp 1694700623
transform 1 0 68208 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_661
timestamp 1694700623
transform 1 0 75376 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_667
timestamp 1694700623
transform 1 0 76048 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_731
timestamp 1694700623
transform 1 0 83216 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_737
timestamp 1694700623
transform 1 0 83888 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_801
timestamp 1694700623
transform 1 0 91056 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_807
timestamp 1694700623
transform 1 0 91728 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_871
timestamp 1694700623
transform 1 0 98896 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_877
timestamp 1694700623
transform 1 0 99568 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_941
timestamp 1694700623
transform 1 0 106736 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_947
timestamp 1694700623
transform 1 0 107408 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1011
timestamp 1694700623
transform 1 0 114576 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1017
timestamp 1694700623
transform 1 0 115248 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1081
timestamp 1694700623
transform 1 0 122416 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1087
timestamp 1694700623
transform 1 0 123088 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1151
timestamp 1694700623
transform 1 0 130256 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1157
timestamp 1694700623
transform 1 0 130928 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1221
timestamp 1694700623
transform 1 0 138096 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1227
timestamp 1694700623
transform 1 0 138768 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1291
timestamp 1694700623
transform 1 0 145936 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1297
timestamp 1694700623
transform 1 0 146608 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1361
timestamp 1694700623
transform 1 0 153776 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1367
timestamp 1694700623
transform 1 0 154448 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1431
timestamp 1694700623
transform 1 0 161616 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1437
timestamp 1694700623
transform 1 0 162288 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1501
timestamp 1694700623
transform 1 0 169456 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1507
timestamp 1694700623
transform 1 0 170128 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1571
timestamp 1694700623
transform 1 0 177296 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1577
timestamp 1694700623
transform 1 0 177968 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1641
timestamp 1694700623
transform 1 0 185136 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1647
timestamp 1694700623
transform 1 0 185808 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1711
timestamp 1694700623
transform 1 0 192976 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_190_1717
timestamp 1694700623
transform 1 0 193648 0 1 152096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_190_1781
timestamp 1694700623
transform 1 0 200816 0 1 152096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_190_1787
timestamp 1694700623
transform 1 0 201488 0 1 152096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_190_1803
timestamp 1694700623
transform 1 0 203280 0 1 152096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190_1811
timestamp 1694700623
transform 1 0 204176 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_190_1813
timestamp 1694700623
transform 1 0 204400 0 1 152096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_2
timestamp 1694700623
transform 1 0 1568 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_66
timestamp 1694700623
transform 1 0 8736 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_72
timestamp 1694700623
transform 1 0 9408 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_136
timestamp 1694700623
transform 1 0 16576 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_142
timestamp 1694700623
transform 1 0 17248 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_206
timestamp 1694700623
transform 1 0 24416 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_212
timestamp 1694700623
transform 1 0 25088 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_276
timestamp 1694700623
transform 1 0 32256 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_282
timestamp 1694700623
transform 1 0 32928 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_346
timestamp 1694700623
transform 1 0 40096 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_352
timestamp 1694700623
transform 1 0 40768 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_416
timestamp 1694700623
transform 1 0 47936 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_422
timestamp 1694700623
transform 1 0 48608 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_486
timestamp 1694700623
transform 1 0 55776 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_492
timestamp 1694700623
transform 1 0 56448 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_556
timestamp 1694700623
transform 1 0 63616 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_562
timestamp 1694700623
transform 1 0 64288 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_626
timestamp 1694700623
transform 1 0 71456 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_632
timestamp 1694700623
transform 1 0 72128 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_696
timestamp 1694700623
transform 1 0 79296 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_702
timestamp 1694700623
transform 1 0 79968 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_766
timestamp 1694700623
transform 1 0 87136 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_772
timestamp 1694700623
transform 1 0 87808 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_836
timestamp 1694700623
transform 1 0 94976 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_842
timestamp 1694700623
transform 1 0 95648 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_906
timestamp 1694700623
transform 1 0 102816 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_912
timestamp 1694700623
transform 1 0 103488 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_976
timestamp 1694700623
transform 1 0 110656 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_982
timestamp 1694700623
transform 1 0 111328 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1046
timestamp 1694700623
transform 1 0 118496 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1052
timestamp 1694700623
transform 1 0 119168 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1116
timestamp 1694700623
transform 1 0 126336 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1122
timestamp 1694700623
transform 1 0 127008 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1186
timestamp 1694700623
transform 1 0 134176 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1192
timestamp 1694700623
transform 1 0 134848 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1256
timestamp 1694700623
transform 1 0 142016 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1262
timestamp 1694700623
transform 1 0 142688 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1326
timestamp 1694700623
transform 1 0 149856 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1332
timestamp 1694700623
transform 1 0 150528 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1396
timestamp 1694700623
transform 1 0 157696 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1402
timestamp 1694700623
transform 1 0 158368 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1466
timestamp 1694700623
transform 1 0 165536 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1472
timestamp 1694700623
transform 1 0 166208 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1536
timestamp 1694700623
transform 1 0 173376 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1542
timestamp 1694700623
transform 1 0 174048 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1606
timestamp 1694700623
transform 1 0 181216 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1612
timestamp 1694700623
transform 1 0 181888 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1676
timestamp 1694700623
transform 1 0 189056 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_191_1682
timestamp 1694700623
transform 1 0 189728 0 -1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1746
timestamp 1694700623
transform 1 0 196896 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_191_1752
timestamp 1694700623
transform 1 0 197568 0 -1 153664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_191_1784
timestamp 1694700623
transform 1 0 201152 0 -1 153664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_191_1800
timestamp 1694700623
transform 1 0 202944 0 -1 153664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_191_1808
timestamp 1694700623
transform 1 0 203840 0 -1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_191_1812
timestamp 1694700623
transform 1 0 204288 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_192_2
timestamp 1694700623
transform 1 0 1568 0 1 153664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192_34
timestamp 1694700623
transform 1 0 5152 0 1 153664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_37
timestamp 1694700623
transform 1 0 5488 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_101
timestamp 1694700623
transform 1 0 12656 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_107
timestamp 1694700623
transform 1 0 13328 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_171
timestamp 1694700623
transform 1 0 20496 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_177
timestamp 1694700623
transform 1 0 21168 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_241
timestamp 1694700623
transform 1 0 28336 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_247
timestamp 1694700623
transform 1 0 29008 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_311
timestamp 1694700623
transform 1 0 36176 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_317
timestamp 1694700623
transform 1 0 36848 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_381
timestamp 1694700623
transform 1 0 44016 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_387
timestamp 1694700623
transform 1 0 44688 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_451
timestamp 1694700623
transform 1 0 51856 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_457
timestamp 1694700623
transform 1 0 52528 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_521
timestamp 1694700623
transform 1 0 59696 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_527
timestamp 1694700623
transform 1 0 60368 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_591
timestamp 1694700623
transform 1 0 67536 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_597
timestamp 1694700623
transform 1 0 68208 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_661
timestamp 1694700623
transform 1 0 75376 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_667
timestamp 1694700623
transform 1 0 76048 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_731
timestamp 1694700623
transform 1 0 83216 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_737
timestamp 1694700623
transform 1 0 83888 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_801
timestamp 1694700623
transform 1 0 91056 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_807
timestamp 1694700623
transform 1 0 91728 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_871
timestamp 1694700623
transform 1 0 98896 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_877
timestamp 1694700623
transform 1 0 99568 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_941
timestamp 1694700623
transform 1 0 106736 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_947
timestamp 1694700623
transform 1 0 107408 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1011
timestamp 1694700623
transform 1 0 114576 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1017
timestamp 1694700623
transform 1 0 115248 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1081
timestamp 1694700623
transform 1 0 122416 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1087
timestamp 1694700623
transform 1 0 123088 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1151
timestamp 1694700623
transform 1 0 130256 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1157
timestamp 1694700623
transform 1 0 130928 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1221
timestamp 1694700623
transform 1 0 138096 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1227
timestamp 1694700623
transform 1 0 138768 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1291
timestamp 1694700623
transform 1 0 145936 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1297
timestamp 1694700623
transform 1 0 146608 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1361
timestamp 1694700623
transform 1 0 153776 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1367
timestamp 1694700623
transform 1 0 154448 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1431
timestamp 1694700623
transform 1 0 161616 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1437
timestamp 1694700623
transform 1 0 162288 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1501
timestamp 1694700623
transform 1 0 169456 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1507
timestamp 1694700623
transform 1 0 170128 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1571
timestamp 1694700623
transform 1 0 177296 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1577
timestamp 1694700623
transform 1 0 177968 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1641
timestamp 1694700623
transform 1 0 185136 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1647
timestamp 1694700623
transform 1 0 185808 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1711
timestamp 1694700623
transform 1 0 192976 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_192_1717
timestamp 1694700623
transform 1 0 193648 0 1 153664
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192_1781
timestamp 1694700623
transform 1 0 200816 0 1 153664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_192_1787
timestamp 1694700623
transform 1 0 201488 0 1 153664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_192_1803
timestamp 1694700623
transform 1 0 203280 0 1 153664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_192_1811
timestamp 1694700623
transform 1 0 204176 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192_1813
timestamp 1694700623
transform 1 0 204400 0 1 153664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_6
timestamp 1694700623
transform 1 0 2016 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_72
timestamp 1694700623
transform 1 0 9408 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_136
timestamp 1694700623
transform 1 0 16576 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_142
timestamp 1694700623
transform 1 0 17248 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_206
timestamp 1694700623
transform 1 0 24416 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_212
timestamp 1694700623
transform 1 0 25088 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_276
timestamp 1694700623
transform 1 0 32256 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_282
timestamp 1694700623
transform 1 0 32928 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_346
timestamp 1694700623
transform 1 0 40096 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_352
timestamp 1694700623
transform 1 0 40768 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_416
timestamp 1694700623
transform 1 0 47936 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_422
timestamp 1694700623
transform 1 0 48608 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_486
timestamp 1694700623
transform 1 0 55776 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_492
timestamp 1694700623
transform 1 0 56448 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_556
timestamp 1694700623
transform 1 0 63616 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_562
timestamp 1694700623
transform 1 0 64288 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_626
timestamp 1694700623
transform 1 0 71456 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_632
timestamp 1694700623
transform 1 0 72128 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_696
timestamp 1694700623
transform 1 0 79296 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_702
timestamp 1694700623
transform 1 0 79968 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_766
timestamp 1694700623
transform 1 0 87136 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_772
timestamp 1694700623
transform 1 0 87808 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_836
timestamp 1694700623
transform 1 0 94976 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_842
timestamp 1694700623
transform 1 0 95648 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_906
timestamp 1694700623
transform 1 0 102816 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_912
timestamp 1694700623
transform 1 0 103488 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_976
timestamp 1694700623
transform 1 0 110656 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_982
timestamp 1694700623
transform 1 0 111328 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1046
timestamp 1694700623
transform 1 0 118496 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1052
timestamp 1694700623
transform 1 0 119168 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1116
timestamp 1694700623
transform 1 0 126336 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1122
timestamp 1694700623
transform 1 0 127008 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1186
timestamp 1694700623
transform 1 0 134176 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1192
timestamp 1694700623
transform 1 0 134848 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1256
timestamp 1694700623
transform 1 0 142016 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1262
timestamp 1694700623
transform 1 0 142688 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1326
timestamp 1694700623
transform 1 0 149856 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1332
timestamp 1694700623
transform 1 0 150528 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1396
timestamp 1694700623
transform 1 0 157696 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1402
timestamp 1694700623
transform 1 0 158368 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1466
timestamp 1694700623
transform 1 0 165536 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1472
timestamp 1694700623
transform 1 0 166208 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1536
timestamp 1694700623
transform 1 0 173376 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1542
timestamp 1694700623
transform 1 0 174048 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1606
timestamp 1694700623
transform 1 0 181216 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1612
timestamp 1694700623
transform 1 0 181888 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1676
timestamp 1694700623
transform 1 0 189056 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_193_1682
timestamp 1694700623
transform 1 0 189728 0 -1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_193_1746
timestamp 1694700623
transform 1 0 196896 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_193_1752
timestamp 1694700623
transform 1 0 197568 0 -1 155232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_193_1784
timestamp 1694700623
transform 1 0 201152 0 -1 155232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_193_1800
timestamp 1694700623
transform 1 0 202944 0 -1 155232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_193_1808
timestamp 1694700623
transform 1 0 203840 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_2
timestamp 1694700623
transform 1 0 1568 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_194_6
timestamp 1694700623
transform 1 0 2016 0 1 155232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_194_22
timestamp 1694700623
transform 1 0 3808 0 1 155232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_30
timestamp 1694700623
transform 1 0 4704 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_194_34
timestamp 1694700623
transform 1 0 5152 0 1 155232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_37
timestamp 1694700623
transform 1 0 5488 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_101
timestamp 1694700623
transform 1 0 12656 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_107
timestamp 1694700623
transform 1 0 13328 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_171
timestamp 1694700623
transform 1 0 20496 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_177
timestamp 1694700623
transform 1 0 21168 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_241
timestamp 1694700623
transform 1 0 28336 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_247
timestamp 1694700623
transform 1 0 29008 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_311
timestamp 1694700623
transform 1 0 36176 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_317
timestamp 1694700623
transform 1 0 36848 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_381
timestamp 1694700623
transform 1 0 44016 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_387
timestamp 1694700623
transform 1 0 44688 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_451
timestamp 1694700623
transform 1 0 51856 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_457
timestamp 1694700623
transform 1 0 52528 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_521
timestamp 1694700623
transform 1 0 59696 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_527
timestamp 1694700623
transform 1 0 60368 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_591
timestamp 1694700623
transform 1 0 67536 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_597
timestamp 1694700623
transform 1 0 68208 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_661
timestamp 1694700623
transform 1 0 75376 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_667
timestamp 1694700623
transform 1 0 76048 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_731
timestamp 1694700623
transform 1 0 83216 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_737
timestamp 1694700623
transform 1 0 83888 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_801
timestamp 1694700623
transform 1 0 91056 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_807
timestamp 1694700623
transform 1 0 91728 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_871
timestamp 1694700623
transform 1 0 98896 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_877
timestamp 1694700623
transform 1 0 99568 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_941
timestamp 1694700623
transform 1 0 106736 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_947
timestamp 1694700623
transform 1 0 107408 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1011
timestamp 1694700623
transform 1 0 114576 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1017
timestamp 1694700623
transform 1 0 115248 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1081
timestamp 1694700623
transform 1 0 122416 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1087
timestamp 1694700623
transform 1 0 123088 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1151
timestamp 1694700623
transform 1 0 130256 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1157
timestamp 1694700623
transform 1 0 130928 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1221
timestamp 1694700623
transform 1 0 138096 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1227
timestamp 1694700623
transform 1 0 138768 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1291
timestamp 1694700623
transform 1 0 145936 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1297
timestamp 1694700623
transform 1 0 146608 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1361
timestamp 1694700623
transform 1 0 153776 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1367
timestamp 1694700623
transform 1 0 154448 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1431
timestamp 1694700623
transform 1 0 161616 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1437
timestamp 1694700623
transform 1 0 162288 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1501
timestamp 1694700623
transform 1 0 169456 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_194_1507
timestamp 1694700623
transform 1 0 170128 0 1 155232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1515
timestamp 1694700623
transform 1 0 171024 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_1545
timestamp 1694700623
transform 1 0 174384 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_194_1549
timestamp 1694700623
transform 1 0 174832 0 1 155232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_194_1565
timestamp 1694700623
transform 1 0 176624 0 1 155232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_1573
timestamp 1694700623
transform 1 0 177520 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1577
timestamp 1694700623
transform 1 0 177968 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1641
timestamp 1694700623
transform 1 0 185136 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_194_1647
timestamp 1694700623
transform 1 0 185808 0 1 155232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1711
timestamp 1694700623
transform 1 0 192976 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_194_1717
timestamp 1694700623
transform 1 0 193648 0 1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_1721
timestamp 1694700623
transform 1 0 194096 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_1749
timestamp 1694700623
transform 1 0 197232 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_194_1753
timestamp 1694700623
transform 1 0 197680 0 1 155232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_194_1787
timestamp 1694700623
transform 1 0 201488 0 1 155232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_194_1803
timestamp 1694700623
transform 1 0 203280 0 1 155232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_194_1811
timestamp 1694700623
transform 1 0 204176 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_194_1813
timestamp 1694700623
transform 1 0 204400 0 1 155232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_16
timestamp 1694700623
transform 1 0 3136 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_20
timestamp 1694700623
transform 1 0 3584 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_22
timestamp 1694700623
transform 1 0 3808 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_27
timestamp 1694700623
transform 1 0 4368 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_31
timestamp 1694700623
transform 1 0 4816 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_33
timestamp 1694700623
transform 1 0 5040 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_36
timestamp 1694700623
transform 1 0 5376 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_70
timestamp 1694700623
transform 1 0 9184 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_86
timestamp 1694700623
transform 1 0 10976 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_90
timestamp 1694700623
transform 1 0 11424 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_95
timestamp 1694700623
transform 1 0 11984 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_99
timestamp 1694700623
transform 1 0 12432 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_101
timestamp 1694700623
transform 1 0 12656 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_104
timestamp 1694700623
transform 1 0 12992 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_138
timestamp 1694700623
transform 1 0 16800 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_154
timestamp 1694700623
transform 1 0 18592 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_156
timestamp 1694700623
transform 1 0 18816 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_169
timestamp 1694700623
transform 1 0 20272 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_172
timestamp 1694700623
transform 1 0 20608 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_206
timestamp 1694700623
transform 1 0 24416 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_222
timestamp 1694700623
transform 1 0 26208 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_226
timestamp 1694700623
transform 1 0 26656 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_231
timestamp 1694700623
transform 1 0 27216 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_235
timestamp 1694700623
transform 1 0 27664 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_237
timestamp 1694700623
transform 1 0 27888 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_240
timestamp 1694700623
transform 1 0 28224 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_274
timestamp 1694700623
transform 1 0 32032 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_290
timestamp 1694700623
transform 1 0 33824 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_294
timestamp 1694700623
transform 1 0 34272 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_299
timestamp 1694700623
transform 1 0 34832 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_303
timestamp 1694700623
transform 1 0 35280 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_305
timestamp 1694700623
transform 1 0 35504 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_308
timestamp 1694700623
transform 1 0 35840 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_342
timestamp 1694700623
transform 1 0 39648 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_358
timestamp 1694700623
transform 1 0 41440 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_376
timestamp 1694700623
transform 1 0 43456 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_380
timestamp 1694700623
transform 1 0 43904 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_396
timestamp 1694700623
transform 1 0 45696 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_404
timestamp 1694700623
transform 1 0 46592 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_410
timestamp 1694700623
transform 1 0 47264 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_426
timestamp 1694700623
transform 1 0 49056 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_430
timestamp 1694700623
transform 1 0 49504 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_435
timestamp 1694700623
transform 1 0 50064 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_439
timestamp 1694700623
transform 1 0 50512 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_441
timestamp 1694700623
transform 1 0 50736 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_444
timestamp 1694700623
transform 1 0 51072 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_478
timestamp 1694700623
transform 1 0 54880 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_494
timestamp 1694700623
transform 1 0 56672 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_498
timestamp 1694700623
transform 1 0 57120 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_503
timestamp 1694700623
transform 1 0 57680 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_507
timestamp 1694700623
transform 1 0 58128 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_509
timestamp 1694700623
transform 1 0 58352 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_512
timestamp 1694700623
transform 1 0 58688 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_546
timestamp 1694700623
transform 1 0 62496 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_562
timestamp 1694700623
transform 1 0 64288 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_580
timestamp 1694700623
transform 1 0 66304 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_584
timestamp 1694700623
transform 1 0 66752 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_600
timestamp 1694700623
transform 1 0 68544 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_608
timestamp 1694700623
transform 1 0 69440 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_614
timestamp 1694700623
transform 1 0 70112 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_630
timestamp 1694700623
transform 1 0 71904 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_634
timestamp 1694700623
transform 1 0 72352 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_639
timestamp 1694700623
transform 1 0 72912 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_643
timestamp 1694700623
transform 1 0 73360 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_645
timestamp 1694700623
transform 1 0 73584 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_648
timestamp 1694700623
transform 1 0 73920 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_682
timestamp 1694700623
transform 1 0 77728 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_698
timestamp 1694700623
transform 1 0 79520 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_702
timestamp 1694700623
transform 1 0 79968 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_707
timestamp 1694700623
transform 1 0 80528 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_711
timestamp 1694700623
transform 1 0 80976 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_713
timestamp 1694700623
transform 1 0 81200 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_716
timestamp 1694700623
transform 1 0 81536 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_750
timestamp 1694700623
transform 1 0 85344 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_766
timestamp 1694700623
transform 1 0 87136 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_784
timestamp 1694700623
transform 1 0 89152 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_788
timestamp 1694700623
transform 1 0 89600 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_804
timestamp 1694700623
transform 1 0 91392 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_812
timestamp 1694700623
transform 1 0 92288 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_818
timestamp 1694700623
transform 1 0 92960 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_834
timestamp 1694700623
transform 1 0 94752 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_838
timestamp 1694700623
transform 1 0 95200 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_843
timestamp 1694700623
transform 1 0 95760 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_847
timestamp 1694700623
transform 1 0 96208 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_849
timestamp 1694700623
transform 1 0 96432 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_852
timestamp 1694700623
transform 1 0 96768 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_886
timestamp 1694700623
transform 1 0 100576 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_902
timestamp 1694700623
transform 1 0 102368 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_906
timestamp 1694700623
transform 1 0 102816 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_911
timestamp 1694700623
transform 1 0 103376 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_915
timestamp 1694700623
transform 1 0 103824 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_917
timestamp 1694700623
transform 1 0 104048 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_920
timestamp 1694700623
transform 1 0 104384 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_954
timestamp 1694700623
transform 1 0 108192 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_970
timestamp 1694700623
transform 1 0 109984 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_972
timestamp 1694700623
transform 1 0 110208 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_985
timestamp 1694700623
transform 1 0 111664 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_988
timestamp 1694700623
transform 1 0 112000 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1022
timestamp 1694700623
transform 1 0 115808 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1038
timestamp 1694700623
transform 1 0 117600 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1042
timestamp 1694700623
transform 1 0 118048 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1047
timestamp 1694700623
transform 1 0 118608 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1051
timestamp 1694700623
transform 1 0 119056 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1053
timestamp 1694700623
transform 1 0 119280 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1056
timestamp 1694700623
transform 1 0 119616 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1090
timestamp 1694700623
transform 1 0 123424 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1106
timestamp 1694700623
transform 1 0 125216 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1110
timestamp 1694700623
transform 1 0 125664 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1115
timestamp 1694700623
transform 1 0 126224 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1119
timestamp 1694700623
transform 1 0 126672 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1121
timestamp 1694700623
transform 1 0 126896 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1124
timestamp 1694700623
transform 1 0 127232 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1158
timestamp 1694700623
transform 1 0 131040 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1174
timestamp 1694700623
transform 1 0 132832 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1192
timestamp 1694700623
transform 1 0 134848 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1196
timestamp 1694700623
transform 1 0 135296 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_1212
timestamp 1694700623
transform 1 0 137088 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1220
timestamp 1694700623
transform 1 0 137984 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1226
timestamp 1694700623
transform 1 0 138656 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1242
timestamp 1694700623
transform 1 0 140448 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1246
timestamp 1694700623
transform 1 0 140896 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1251
timestamp 1694700623
transform 1 0 141456 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1255
timestamp 1694700623
transform 1 0 141904 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1257
timestamp 1694700623
transform 1 0 142128 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1260
timestamp 1694700623
transform 1 0 142464 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1294
timestamp 1694700623
transform 1 0 146272 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1310
timestamp 1694700623
transform 1 0 148064 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1314
timestamp 1694700623
transform 1 0 148512 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1319
timestamp 1694700623
transform 1 0 149072 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1323
timestamp 1694700623
transform 1 0 149520 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1325
timestamp 1694700623
transform 1 0 149744 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1328
timestamp 1694700623
transform 1 0 150080 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1362
timestamp 1694700623
transform 1 0 153888 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1378
timestamp 1694700623
transform 1 0 155680 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1396
timestamp 1694700623
transform 1 0 157696 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1400
timestamp 1694700623
transform 1 0 158144 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_1416
timestamp 1694700623
transform 1 0 159936 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1424
timestamp 1694700623
transform 1 0 160832 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1430
timestamp 1694700623
transform 1 0 161504 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1446
timestamp 1694700623
transform 1 0 163296 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1450
timestamp 1694700623
transform 1 0 163744 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1455
timestamp 1694700623
transform 1 0 164304 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1459
timestamp 1694700623
transform 1 0 164752 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1461
timestamp 1694700623
transform 1 0 164976 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1464
timestamp 1694700623
transform 1 0 165312 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1498
timestamp 1694700623
transform 1 0 169120 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1532
timestamp 1694700623
transform 1 0 172928 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1566
timestamp 1694700623
transform 1 0 176736 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1600
timestamp 1694700623
transform 1 0 180544 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_195_1634
timestamp 1694700623
transform 1 0 184352 0 -1 156800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1650
timestamp 1694700623
transform 1 0 186144 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1654
timestamp 1694700623
transform 1 0 186592 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_195_1659
timestamp 1694700623
transform 1 0 187152 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1663
timestamp 1694700623
transform 1 0 187600 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_195_1665
timestamp 1694700623
transform 1 0 187824 0 -1 156800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1668
timestamp 1694700623
transform 1 0 188160 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1702
timestamp 1694700623
transform 1 0 191968 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1736
timestamp 1694700623
transform 1 0 195776 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_195_1770
timestamp 1694700623
transform 1 0 199584 0 -1 156800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195_1804
timestamp 1694700623
transform 1 0 203392 0 -1 156800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195_1812
timestamp 1694700623
transform 1 0 204288 0 -1 156800
box -86 -86 310 870
use gf180_sram_8x1024  gf180_sram_8x1024
timestamp 0
transform 1 0 20000 0 1 20000
box 0 0 166264 122572
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input1 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 110544 0 -1 156800
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input2 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 88928 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input3
timestamp 1694700623
transform 1 0 64512 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  input4 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 41664 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input5
timestamp 1694700623
transform 1 0 19152 0 -1 156800
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input6 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input7
timestamp 1694700623
transform 1 0 1568 0 -1 147392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input8
timestamp 1694700623
transform 1 0 1568 0 1 134848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input9
timestamp 1694700623
transform 1 0 1568 0 1 123872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input10
timestamp 1694700623
transform 1 0 1568 0 -1 112896
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 101920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1694700623
transform 1 0 1568 0 1 89376
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1694700623
transform 1 0 1568 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1694700623
transform 1 0 1568 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1694700623
transform 1 0 1568 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1694700623
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1694700623
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input20
timestamp 1694700623
transform -1 0 157472 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input21
timestamp 1694700623
transform -1 0 134624 0 -1 156800
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 201600 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1694700623
transform 1 0 201600 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1694700623
transform 1 0 201040 0 -1 67424
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1694700623
transform 1 0 201040 0 -1 94080
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1694700623
transform 1 0 201600 0 1 119168
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1694700623
transform 1 0 201600 0 1 145824
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1694700623
transform -1 0 197232 0 1 155232
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1694700623
transform -1 0 174384 0 1 155232
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_196 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 204736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_197
timestamp 1694700623
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 204736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_198
timestamp 1694700623
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 204736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_199
timestamp 1694700623
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 204736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_200
timestamp 1694700623
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 204736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_201
timestamp 1694700623
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 204736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_202
timestamp 1694700623
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 204736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_203
timestamp 1694700623
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 204736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_204
timestamp 1694700623
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 204736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_205
timestamp 1694700623
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 204736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_206
timestamp 1694700623
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 204736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_207
timestamp 1694700623
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 204736 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_208
timestamp 1694700623
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 204736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_209
timestamp 1694700623
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 204736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_210
timestamp 1694700623
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 204736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_211
timestamp 1694700623
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 204736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_212
timestamp 1694700623
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 204736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_213
timestamp 1694700623
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 204736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_1_Left_391
timestamp 1694700623
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_1_Right_717
timestamp 1694700623
transform -1 0 17920 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_2_Left_392
timestamp 1694700623
transform 1 0 188272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_2_Right_33
timestamp 1694700623
transform -1 0 204736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_1_Left_214
timestamp 1694700623
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_1_Right_555
timestamp 1694700623
transform -1 0 17920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_2_Left_393
timestamp 1694700623
transform 1 0 188272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_2_Right_34
timestamp 1694700623
transform -1 0 204736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_1_Left_215
timestamp 1694700623
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_1_Right_556
timestamp 1694700623
transform -1 0 17920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_2_Left_394
timestamp 1694700623
transform 1 0 188272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_2_Right_35
timestamp 1694700623
transform -1 0 204736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_1_Left_216
timestamp 1694700623
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_1_Right_557
timestamp 1694700623
transform -1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_2_Left_395
timestamp 1694700623
transform 1 0 188272 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_2_Right_36
timestamp 1694700623
transform -1 0 204736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_1_Left_217
timestamp 1694700623
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_1_Right_558
timestamp 1694700623
transform -1 0 17920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_2_Left_396
timestamp 1694700623
transform 1 0 188272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_2_Right_37
timestamp 1694700623
transform -1 0 204736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_1_Left_218
timestamp 1694700623
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_1_Right_559
timestamp 1694700623
transform -1 0 17920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_2_Left_397
timestamp 1694700623
transform 1 0 188272 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_2_Right_38
timestamp 1694700623
transform -1 0 204736 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_1_Left_219
timestamp 1694700623
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_1_Right_560
timestamp 1694700623
transform -1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_2_Left_398
timestamp 1694700623
transform 1 0 188272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_2_Right_39
timestamp 1694700623
transform -1 0 204736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_1_Left_220
timestamp 1694700623
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_1_Right_561
timestamp 1694700623
transform -1 0 17920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_2_Left_399
timestamp 1694700623
transform 1 0 188272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_2_Right_40
timestamp 1694700623
transform -1 0 204736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_1_Left_221
timestamp 1694700623
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_1_Right_562
timestamp 1694700623
transform -1 0 17920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_2_Left_400
timestamp 1694700623
transform 1 0 188272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_2_Right_41
timestamp 1694700623
transform -1 0 204736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_1_Left_222
timestamp 1694700623
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_1_Right_563
timestamp 1694700623
transform -1 0 17920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_2_Left_401
timestamp 1694700623
transform 1 0 188272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_2_Right_42
timestamp 1694700623
transform -1 0 204736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_1_Left_223
timestamp 1694700623
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_1_Right_564
timestamp 1694700623
transform -1 0 17920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_2_Left_402
timestamp 1694700623
transform 1 0 188272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_2_Right_43
timestamp 1694700623
transform -1 0 204736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_1_Left_224
timestamp 1694700623
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_1_Right_565
timestamp 1694700623
transform -1 0 17920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_2_Left_403
timestamp 1694700623
transform 1 0 188272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_2_Right_44
timestamp 1694700623
transform -1 0 204736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_1_Left_225
timestamp 1694700623
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_1_Right_566
timestamp 1694700623
transform -1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_2_Left_404
timestamp 1694700623
transform 1 0 188272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_2_Right_45
timestamp 1694700623
transform -1 0 204736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_1_Left_226
timestamp 1694700623
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_1_Right_567
timestamp 1694700623
transform -1 0 17920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_2_Left_405
timestamp 1694700623
transform 1 0 188272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_2_Right_46
timestamp 1694700623
transform -1 0 204736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_1_Left_227
timestamp 1694700623
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_1_Right_568
timestamp 1694700623
transform -1 0 17920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_2_Left_406
timestamp 1694700623
transform 1 0 188272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_2_Right_47
timestamp 1694700623
transform -1 0 204736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_1_Left_228
timestamp 1694700623
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_1_Right_569
timestamp 1694700623
transform -1 0 17920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_2_Left_407
timestamp 1694700623
transform 1 0 188272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_2_Right_48
timestamp 1694700623
transform -1 0 204736 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_1_Left_229
timestamp 1694700623
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_1_Right_570
timestamp 1694700623
transform -1 0 17920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_2_Left_408
timestamp 1694700623
transform 1 0 188272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_2_Right_49
timestamp 1694700623
transform -1 0 204736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_1_Left_230
timestamp 1694700623
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_1_Right_571
timestamp 1694700623
transform -1 0 17920 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_2_Left_409
timestamp 1694700623
transform 1 0 188272 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_2_Right_50
timestamp 1694700623
transform -1 0 204736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_1_Left_231
timestamp 1694700623
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_1_Right_572
timestamp 1694700623
transform -1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_2_Left_410
timestamp 1694700623
transform 1 0 188272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_2_Right_51
timestamp 1694700623
transform -1 0 204736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_1_Left_232
timestamp 1694700623
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_1_Right_573
timestamp 1694700623
transform -1 0 17920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_2_Left_411
timestamp 1694700623
transform 1 0 188272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_2_Right_52
timestamp 1694700623
transform -1 0 204736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_1_Left_233
timestamp 1694700623
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_1_Right_574
timestamp 1694700623
transform -1 0 17920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_2_Left_412
timestamp 1694700623
transform 1 0 188272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_2_Right_53
timestamp 1694700623
transform -1 0 204736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_1_Left_234
timestamp 1694700623
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_1_Right_575
timestamp 1694700623
transform -1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_2_Left_413
timestamp 1694700623
transform 1 0 188272 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_2_Right_54
timestamp 1694700623
transform -1 0 204736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_1_Left_235
timestamp 1694700623
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_1_Right_576
timestamp 1694700623
transform -1 0 17920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_2_Left_414
timestamp 1694700623
transform 1 0 188272 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_2_Right_55
timestamp 1694700623
transform -1 0 204736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_1_Left_236
timestamp 1694700623
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_1_Right_577
timestamp 1694700623
transform -1 0 17920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_2_Left_415
timestamp 1694700623
transform 1 0 188272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_2_Right_56
timestamp 1694700623
transform -1 0 204736 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_1_Left_237
timestamp 1694700623
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_1_Right_578
timestamp 1694700623
transform -1 0 17920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_2_Left_416
timestamp 1694700623
transform 1 0 188272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_2_Right_57
timestamp 1694700623
transform -1 0 204736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_1_Left_238
timestamp 1694700623
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_1_Right_579
timestamp 1694700623
transform -1 0 17920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_2_Left_417
timestamp 1694700623
transform 1 0 188272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_2_Right_58
timestamp 1694700623
transform -1 0 204736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_1_Left_239
timestamp 1694700623
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_1_Right_580
timestamp 1694700623
transform -1 0 17920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_2_Left_418
timestamp 1694700623
transform 1 0 188272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_2_Right_59
timestamp 1694700623
transform -1 0 204736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_1_Left_240
timestamp 1694700623
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_1_Right_581
timestamp 1694700623
transform -1 0 17920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_2_Left_419
timestamp 1694700623
transform 1 0 188272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_2_Right_60
timestamp 1694700623
transform -1 0 204736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_1_Left_241
timestamp 1694700623
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_1_Right_582
timestamp 1694700623
transform -1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_2_Left_420
timestamp 1694700623
transform 1 0 188272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_2_Right_61
timestamp 1694700623
transform -1 0 204736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_1_Left_242
timestamp 1694700623
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_1_Right_583
timestamp 1694700623
transform -1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_2_Left_421
timestamp 1694700623
transform 1 0 188272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_2_Right_62
timestamp 1694700623
transform -1 0 204736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_1_Left_243
timestamp 1694700623
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_1_Right_584
timestamp 1694700623
transform -1 0 17920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_2_Left_422
timestamp 1694700623
transform 1 0 188272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_2_Right_63
timestamp 1694700623
transform -1 0 204736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_1_Left_244
timestamp 1694700623
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_1_Right_585
timestamp 1694700623
transform -1 0 17920 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_2_Left_423
timestamp 1694700623
transform 1 0 188272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_2_Right_64
timestamp 1694700623
transform -1 0 204736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_1_Left_245
timestamp 1694700623
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_1_Right_586
timestamp 1694700623
transform -1 0 17920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_2_Left_424
timestamp 1694700623
transform 1 0 188272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_2_Right_65
timestamp 1694700623
transform -1 0 204736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_1_Left_246
timestamp 1694700623
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_1_Right_587
timestamp 1694700623
transform -1 0 17920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_2_Left_425
timestamp 1694700623
transform 1 0 188272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_2_Right_66
timestamp 1694700623
transform -1 0 204736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_1_Left_247
timestamp 1694700623
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_1_Right_588
timestamp 1694700623
transform -1 0 17920 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_2_Left_426
timestamp 1694700623
transform 1 0 188272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_2_Right_67
timestamp 1694700623
transform -1 0 204736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_1_Left_248
timestamp 1694700623
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_1_Right_589
timestamp 1694700623
transform -1 0 17920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_2_Left_427
timestamp 1694700623
transform 1 0 188272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_2_Right_68
timestamp 1694700623
transform -1 0 204736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_1_Left_249
timestamp 1694700623
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_1_Right_590
timestamp 1694700623
transform -1 0 17920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_2_Left_428
timestamp 1694700623
transform 1 0 188272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_2_Right_69
timestamp 1694700623
transform -1 0 204736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_1_Left_250
timestamp 1694700623
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_1_Right_591
timestamp 1694700623
transform -1 0 17920 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_2_Left_429
timestamp 1694700623
transform 1 0 188272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_2_Right_70
timestamp 1694700623
transform -1 0 204736 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_1_Left_251
timestamp 1694700623
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_1_Right_592
timestamp 1694700623
transform -1 0 17920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_2_Left_430
timestamp 1694700623
transform 1 0 188272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_2_Right_71
timestamp 1694700623
transform -1 0 204736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_1_Left_252
timestamp 1694700623
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_1_Right_593
timestamp 1694700623
transform -1 0 17920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_2_Left_431
timestamp 1694700623
transform 1 0 188272 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_2_Right_72
timestamp 1694700623
transform -1 0 204736 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_1_Left_253
timestamp 1694700623
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_1_Right_594
timestamp 1694700623
transform -1 0 17920 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_2_Left_432
timestamp 1694700623
transform 1 0 188272 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_2_Right_73
timestamp 1694700623
transform -1 0 204736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_1_Left_254
timestamp 1694700623
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_1_Right_595
timestamp 1694700623
transform -1 0 17920 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_2_Left_433
timestamp 1694700623
transform 1 0 188272 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_2_Right_74
timestamp 1694700623
transform -1 0 204736 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_1_Left_255
timestamp 1694700623
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_1_Right_596
timestamp 1694700623
transform -1 0 17920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_2_Left_434
timestamp 1694700623
transform 1 0 188272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_2_Right_75
timestamp 1694700623
transform -1 0 204736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_1_Left_256
timestamp 1694700623
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_1_Right_597
timestamp 1694700623
transform -1 0 17920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_2_Left_435
timestamp 1694700623
transform 1 0 188272 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_2_Right_76
timestamp 1694700623
transform -1 0 204736 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_1_Left_257
timestamp 1694700623
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_1_Right_598
timestamp 1694700623
transform -1 0 17920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_2_Left_436
timestamp 1694700623
transform 1 0 188272 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_2_Right_77
timestamp 1694700623
transform -1 0 204736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_1_Left_258
timestamp 1694700623
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_1_Right_599
timestamp 1694700623
transform -1 0 17920 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_2_Left_437
timestamp 1694700623
transform 1 0 188272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_2_Right_78
timestamp 1694700623
transform -1 0 204736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_1_Left_259
timestamp 1694700623
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_1_Right_600
timestamp 1694700623
transform -1 0 17920 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_2_Left_438
timestamp 1694700623
transform 1 0 188272 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_2_Right_79
timestamp 1694700623
transform -1 0 204736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_1_Left_260
timestamp 1694700623
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_1_Right_601
timestamp 1694700623
transform -1 0 17920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_2_Left_439
timestamp 1694700623
transform 1 0 188272 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_2_Right_80
timestamp 1694700623
transform -1 0 204736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_1_Left_261
timestamp 1694700623
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_1_Right_602
timestamp 1694700623
transform -1 0 17920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_2_Left_440
timestamp 1694700623
transform 1 0 188272 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_2_Right_81
timestamp 1694700623
transform -1 0 204736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_1_Left_262
timestamp 1694700623
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_1_Right_603
timestamp 1694700623
transform -1 0 17920 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_2_Left_441
timestamp 1694700623
transform 1 0 188272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_2_Right_82
timestamp 1694700623
transform -1 0 204736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_1_Left_263
timestamp 1694700623
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_1_Right_604
timestamp 1694700623
transform -1 0 17920 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_2_Left_442
timestamp 1694700623
transform 1 0 188272 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_2_Right_83
timestamp 1694700623
transform -1 0 204736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_1_Left_264
timestamp 1694700623
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_1_Right_605
timestamp 1694700623
transform -1 0 17920 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_2_Left_443
timestamp 1694700623
transform 1 0 188272 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_2_Right_84
timestamp 1694700623
transform -1 0 204736 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_1_Left_265
timestamp 1694700623
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_1_Right_606
timestamp 1694700623
transform -1 0 17920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_2_Left_444
timestamp 1694700623
transform 1 0 188272 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_2_Right_85
timestamp 1694700623
transform -1 0 204736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_1_Left_266
timestamp 1694700623
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_1_Right_607
timestamp 1694700623
transform -1 0 17920 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_2_Left_445
timestamp 1694700623
transform 1 0 188272 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_2_Right_86
timestamp 1694700623
transform -1 0 204736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_1_Left_267
timestamp 1694700623
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_1_Right_608
timestamp 1694700623
transform -1 0 17920 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_2_Left_446
timestamp 1694700623
transform 1 0 188272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_2_Right_87
timestamp 1694700623
transform -1 0 204736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_1_Left_268
timestamp 1694700623
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_1_Right_609
timestamp 1694700623
transform -1 0 17920 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_2_Left_447
timestamp 1694700623
transform 1 0 188272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_2_Right_88
timestamp 1694700623
transform -1 0 204736 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_1_Left_269
timestamp 1694700623
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_1_Right_610
timestamp 1694700623
transform -1 0 17920 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_2_Left_448
timestamp 1694700623
transform 1 0 188272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_2_Right_89
timestamp 1694700623
transform -1 0 204736 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_1_Left_270
timestamp 1694700623
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_1_Right_611
timestamp 1694700623
transform -1 0 17920 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_2_Left_449
timestamp 1694700623
transform 1 0 188272 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_2_Right_90
timestamp 1694700623
transform -1 0 204736 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_1_Left_271
timestamp 1694700623
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_1_Right_612
timestamp 1694700623
transform -1 0 17920 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_2_Left_450
timestamp 1694700623
transform 1 0 188272 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_2_Right_91
timestamp 1694700623
transform -1 0 204736 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_1_Left_272
timestamp 1694700623
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_1_Right_613
timestamp 1694700623
transform -1 0 17920 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_2_Left_451
timestamp 1694700623
transform 1 0 188272 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_2_Right_92
timestamp 1694700623
transform -1 0 204736 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_1_Left_273
timestamp 1694700623
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_1_Right_614
timestamp 1694700623
transform -1 0 17920 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_2_Left_452
timestamp 1694700623
transform 1 0 188272 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_2_Right_93
timestamp 1694700623
transform -1 0 204736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_1_Left_274
timestamp 1694700623
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_1_Right_615
timestamp 1694700623
transform -1 0 17920 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_2_Left_453
timestamp 1694700623
transform 1 0 188272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_2_Right_94
timestamp 1694700623
transform -1 0 204736 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_1_Left_275
timestamp 1694700623
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_1_Right_616
timestamp 1694700623
transform -1 0 17920 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_2_Left_454
timestamp 1694700623
transform 1 0 188272 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_2_Right_95
timestamp 1694700623
transform -1 0 204736 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_1_Left_276
timestamp 1694700623
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_1_Right_617
timestamp 1694700623
transform -1 0 17920 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_2_Left_455
timestamp 1694700623
transform 1 0 188272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_2_Right_96
timestamp 1694700623
transform -1 0 204736 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_1_Left_277
timestamp 1694700623
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_1_Right_618
timestamp 1694700623
transform -1 0 17920 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_2_Left_456
timestamp 1694700623
transform 1 0 188272 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_2_Right_97
timestamp 1694700623
transform -1 0 204736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_1_Left_278
timestamp 1694700623
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_1_Right_619
timestamp 1694700623
transform -1 0 17920 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_2_Left_457
timestamp 1694700623
transform 1 0 188272 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_2_Right_98
timestamp 1694700623
transform -1 0 204736 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_1_Left_279
timestamp 1694700623
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_1_Right_620
timestamp 1694700623
transform -1 0 17920 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_2_Left_458
timestamp 1694700623
transform 1 0 188272 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_2_Right_99
timestamp 1694700623
transform -1 0 204736 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_1_Left_280
timestamp 1694700623
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_1_Right_621
timestamp 1694700623
transform -1 0 17920 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_2_Left_459
timestamp 1694700623
transform 1 0 188272 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_2_Right_100
timestamp 1694700623
transform -1 0 204736 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_1_Left_281
timestamp 1694700623
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_1_Right_622
timestamp 1694700623
transform -1 0 17920 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_2_Left_460
timestamp 1694700623
transform 1 0 188272 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_2_Right_101
timestamp 1694700623
transform -1 0 204736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_1_Left_282
timestamp 1694700623
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_1_Right_623
timestamp 1694700623
transform -1 0 17920 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_2_Left_461
timestamp 1694700623
transform 1 0 188272 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_2_Right_102
timestamp 1694700623
transform -1 0 204736 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_1_Left_283
timestamp 1694700623
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_1_Right_624
timestamp 1694700623
transform -1 0 17920 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_2_Left_462
timestamp 1694700623
transform 1 0 188272 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_2_Right_103
timestamp 1694700623
transform -1 0 204736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_1_Left_284
timestamp 1694700623
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_1_Right_625
timestamp 1694700623
transform -1 0 17920 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_2_Left_463
timestamp 1694700623
transform 1 0 188272 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_2_Right_104
timestamp 1694700623
transform -1 0 204736 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_1_Left_285
timestamp 1694700623
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_1_Right_626
timestamp 1694700623
transform -1 0 17920 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_2_Left_464
timestamp 1694700623
transform 1 0 188272 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_2_Right_105
timestamp 1694700623
transform -1 0 204736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_1_Left_286
timestamp 1694700623
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_1_Right_627
timestamp 1694700623
transform -1 0 17920 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_2_Left_465
timestamp 1694700623
transform 1 0 188272 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_2_Right_106
timestamp 1694700623
transform -1 0 204736 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_1_Left_287
timestamp 1694700623
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_1_Right_628
timestamp 1694700623
transform -1 0 17920 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_2_Left_466
timestamp 1694700623
transform 1 0 188272 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_2_Right_107
timestamp 1694700623
transform -1 0 204736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_1_Left_288
timestamp 1694700623
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_1_Right_629
timestamp 1694700623
transform -1 0 17920 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_2_Left_467
timestamp 1694700623
transform 1 0 188272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_2_Right_108
timestamp 1694700623
transform -1 0 204736 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_1_Left_289
timestamp 1694700623
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_1_Right_630
timestamp 1694700623
transform -1 0 17920 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_2_Left_468
timestamp 1694700623
transform 1 0 188272 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_2_Right_109
timestamp 1694700623
transform -1 0 204736 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_1_Left_290
timestamp 1694700623
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_1_Right_631
timestamp 1694700623
transform -1 0 17920 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_2_Left_469
timestamp 1694700623
transform 1 0 188272 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_2_Right_110
timestamp 1694700623
transform -1 0 204736 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_1_Left_291
timestamp 1694700623
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_1_Right_632
timestamp 1694700623
transform -1 0 17920 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_2_Left_470
timestamp 1694700623
transform 1 0 188272 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_2_Right_111
timestamp 1694700623
transform -1 0 204736 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_1_Left_292
timestamp 1694700623
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_1_Right_633
timestamp 1694700623
transform -1 0 17920 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_2_Left_471
timestamp 1694700623
transform 1 0 188272 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_2_Right_112
timestamp 1694700623
transform -1 0 204736 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_1_Left_293
timestamp 1694700623
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_1_Right_634
timestamp 1694700623
transform -1 0 17920 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_2_Left_472
timestamp 1694700623
transform 1 0 188272 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_2_Right_113
timestamp 1694700623
transform -1 0 204736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_1_Left_294
timestamp 1694700623
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_1_Right_635
timestamp 1694700623
transform -1 0 17920 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_2_Left_473
timestamp 1694700623
transform 1 0 188272 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_2_Right_114
timestamp 1694700623
transform -1 0 204736 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_1_Left_295
timestamp 1694700623
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_1_Right_636
timestamp 1694700623
transform -1 0 17920 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_2_Left_474
timestamp 1694700623
transform 1 0 188272 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_2_Right_115
timestamp 1694700623
transform -1 0 204736 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_1_Left_296
timestamp 1694700623
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_1_Right_637
timestamp 1694700623
transform -1 0 17920 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_2_Left_475
timestamp 1694700623
transform 1 0 188272 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_2_Right_116
timestamp 1694700623
transform -1 0 204736 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_1_Left_297
timestamp 1694700623
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_1_Right_638
timestamp 1694700623
transform -1 0 17920 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_2_Left_476
timestamp 1694700623
transform 1 0 188272 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_2_Right_117
timestamp 1694700623
transform -1 0 204736 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_1_Left_298
timestamp 1694700623
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_1_Right_639
timestamp 1694700623
transform -1 0 17920 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_2_Left_477
timestamp 1694700623
transform 1 0 188272 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_2_Right_118
timestamp 1694700623
transform -1 0 204736 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_1_Left_299
timestamp 1694700623
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_1_Right_640
timestamp 1694700623
transform -1 0 17920 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_2_Left_478
timestamp 1694700623
transform 1 0 188272 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_2_Right_119
timestamp 1694700623
transform -1 0 204736 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_1_Left_300
timestamp 1694700623
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_1_Right_641
timestamp 1694700623
transform -1 0 17920 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_2_Left_479
timestamp 1694700623
transform 1 0 188272 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_2_Right_120
timestamp 1694700623
transform -1 0 204736 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_1_Left_301
timestamp 1694700623
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_1_Right_642
timestamp 1694700623
transform -1 0 17920 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_2_Left_480
timestamp 1694700623
transform 1 0 188272 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_2_Right_121
timestamp 1694700623
transform -1 0 204736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_1_Left_302
timestamp 1694700623
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_1_Right_643
timestamp 1694700623
transform -1 0 17920 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_2_Left_481
timestamp 1694700623
transform 1 0 188272 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_2_Right_122
timestamp 1694700623
transform -1 0 204736 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_1_Left_303
timestamp 1694700623
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_1_Right_644
timestamp 1694700623
transform -1 0 17920 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_2_Left_482
timestamp 1694700623
transform 1 0 188272 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_2_Right_123
timestamp 1694700623
transform -1 0 204736 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_1_Left_304
timestamp 1694700623
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_1_Right_645
timestamp 1694700623
transform -1 0 17920 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_2_Left_483
timestamp 1694700623
transform 1 0 188272 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_2_Right_124
timestamp 1694700623
transform -1 0 204736 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_1_Left_305
timestamp 1694700623
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_1_Right_646
timestamp 1694700623
transform -1 0 17920 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_2_Left_484
timestamp 1694700623
transform 1 0 188272 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_2_Right_125
timestamp 1694700623
transform -1 0 204736 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_1_Left_306
timestamp 1694700623
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_1_Right_647
timestamp 1694700623
transform -1 0 17920 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_2_Left_485
timestamp 1694700623
transform 1 0 188272 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_2_Right_126
timestamp 1694700623
transform -1 0 204736 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_1_Left_307
timestamp 1694700623
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_1_Right_648
timestamp 1694700623
transform -1 0 17920 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_2_Left_486
timestamp 1694700623
transform 1 0 188272 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_2_Right_127
timestamp 1694700623
transform -1 0 204736 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_1_Left_308
timestamp 1694700623
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_1_Right_649
timestamp 1694700623
transform -1 0 17920 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_2_Left_487
timestamp 1694700623
transform 1 0 188272 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_2_Right_128
timestamp 1694700623
transform -1 0 204736 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_1_Left_309
timestamp 1694700623
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_1_Right_650
timestamp 1694700623
transform -1 0 17920 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_2_Left_488
timestamp 1694700623
transform 1 0 188272 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_2_Right_129
timestamp 1694700623
transform -1 0 204736 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_1_Left_310
timestamp 1694700623
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_1_Right_651
timestamp 1694700623
transform -1 0 17920 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_2_Left_489
timestamp 1694700623
transform 1 0 188272 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_2_Right_130
timestamp 1694700623
transform -1 0 204736 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_1_Left_311
timestamp 1694700623
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_1_Right_652
timestamp 1694700623
transform -1 0 17920 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_2_Left_490
timestamp 1694700623
transform 1 0 188272 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_2_Right_131
timestamp 1694700623
transform -1 0 204736 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_1_Left_312
timestamp 1694700623
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_1_Right_653
timestamp 1694700623
transform -1 0 17920 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_2_Left_491
timestamp 1694700623
transform 1 0 188272 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_2_Right_132
timestamp 1694700623
transform -1 0 204736 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_1_Left_313
timestamp 1694700623
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_1_Right_654
timestamp 1694700623
transform -1 0 17920 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_2_Left_492
timestamp 1694700623
transform 1 0 188272 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_2_Right_133
timestamp 1694700623
transform -1 0 204736 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_1_Left_314
timestamp 1694700623
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_1_Right_655
timestamp 1694700623
transform -1 0 17920 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_2_Left_493
timestamp 1694700623
transform 1 0 188272 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_2_Right_134
timestamp 1694700623
transform -1 0 204736 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_1_Left_315
timestamp 1694700623
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_1_Right_656
timestamp 1694700623
transform -1 0 17920 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_2_Left_494
timestamp 1694700623
transform 1 0 188272 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_2_Right_135
timestamp 1694700623
transform -1 0 204736 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_1_Left_316
timestamp 1694700623
transform 1 0 1344 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_1_Right_657
timestamp 1694700623
transform -1 0 17920 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_2_Left_495
timestamp 1694700623
transform 1 0 188272 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_2_Right_136
timestamp 1694700623
transform -1 0 204736 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_1_Left_317
timestamp 1694700623
transform 1 0 1344 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_1_Right_658
timestamp 1694700623
transform -1 0 17920 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_2_Left_496
timestamp 1694700623
transform 1 0 188272 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_2_Right_137
timestamp 1694700623
transform -1 0 204736 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_1_Left_318
timestamp 1694700623
transform 1 0 1344 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_1_Right_659
timestamp 1694700623
transform -1 0 17920 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_2_Left_497
timestamp 1694700623
transform 1 0 188272 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_2_Right_138
timestamp 1694700623
transform -1 0 204736 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_1_Left_319
timestamp 1694700623
transform 1 0 1344 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_1_Right_660
timestamp 1694700623
transform -1 0 17920 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_2_Left_498
timestamp 1694700623
transform 1 0 188272 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_2_Right_139
timestamp 1694700623
transform -1 0 204736 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_1_Left_320
timestamp 1694700623
transform 1 0 1344 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_1_Right_661
timestamp 1694700623
transform -1 0 17920 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_2_Left_499
timestamp 1694700623
transform 1 0 188272 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_2_Right_140
timestamp 1694700623
transform -1 0 204736 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_1_Left_321
timestamp 1694700623
transform 1 0 1344 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_1_Right_662
timestamp 1694700623
transform -1 0 17920 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_2_Left_500
timestamp 1694700623
transform 1 0 188272 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_2_Right_141
timestamp 1694700623
transform -1 0 204736 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_1_Left_322
timestamp 1694700623
transform 1 0 1344 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_1_Right_663
timestamp 1694700623
transform -1 0 17920 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_2_Left_501
timestamp 1694700623
transform 1 0 188272 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_2_Right_142
timestamp 1694700623
transform -1 0 204736 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_1_Left_323
timestamp 1694700623
transform 1 0 1344 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_1_Right_664
timestamp 1694700623
transform -1 0 17920 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_2_Left_502
timestamp 1694700623
transform 1 0 188272 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_2_Right_143
timestamp 1694700623
transform -1 0 204736 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_1_Left_324
timestamp 1694700623
transform 1 0 1344 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_1_Right_665
timestamp 1694700623
transform -1 0 17920 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_2_Left_503
timestamp 1694700623
transform 1 0 188272 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_2_Right_144
timestamp 1694700623
transform -1 0 204736 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_1_Left_325
timestamp 1694700623
transform 1 0 1344 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_1_Right_666
timestamp 1694700623
transform -1 0 17920 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_2_Left_504
timestamp 1694700623
transform 1 0 188272 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_2_Right_145
timestamp 1694700623
transform -1 0 204736 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_1_Left_326
timestamp 1694700623
transform 1 0 1344 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_1_Right_667
timestamp 1694700623
transform -1 0 17920 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_2_Left_505
timestamp 1694700623
transform 1 0 188272 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_2_Right_146
timestamp 1694700623
transform -1 0 204736 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_1_Left_327
timestamp 1694700623
transform 1 0 1344 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_1_Right_668
timestamp 1694700623
transform -1 0 17920 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_2_Left_506
timestamp 1694700623
transform 1 0 188272 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_2_Right_147
timestamp 1694700623
transform -1 0 204736 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_1_Left_328
timestamp 1694700623
transform 1 0 1344 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_1_Right_669
timestamp 1694700623
transform -1 0 17920 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_2_Left_507
timestamp 1694700623
transform 1 0 188272 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_2_Right_148
timestamp 1694700623
transform -1 0 204736 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_1_Left_329
timestamp 1694700623
transform 1 0 1344 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_1_Right_670
timestamp 1694700623
transform -1 0 17920 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_2_Left_508
timestamp 1694700623
transform 1 0 188272 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_2_Right_149
timestamp 1694700623
transform -1 0 204736 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_1_Left_330
timestamp 1694700623
transform 1 0 1344 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_1_Right_671
timestamp 1694700623
transform -1 0 17920 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_2_Left_509
timestamp 1694700623
transform 1 0 188272 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_2_Right_150
timestamp 1694700623
transform -1 0 204736 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_1_Left_331
timestamp 1694700623
transform 1 0 1344 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_1_Right_672
timestamp 1694700623
transform -1 0 17920 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_2_Left_510
timestamp 1694700623
transform 1 0 188272 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_2_Right_151
timestamp 1694700623
transform -1 0 204736 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_1_Left_332
timestamp 1694700623
transform 1 0 1344 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_1_Right_673
timestamp 1694700623
transform -1 0 17920 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_2_Left_511
timestamp 1694700623
transform 1 0 188272 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_2_Right_152
timestamp 1694700623
transform -1 0 204736 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_1_Left_333
timestamp 1694700623
transform 1 0 1344 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_1_Right_674
timestamp 1694700623
transform -1 0 17920 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_2_Left_512
timestamp 1694700623
transform 1 0 188272 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_2_Right_153
timestamp 1694700623
transform -1 0 204736 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_1_Left_334
timestamp 1694700623
transform 1 0 1344 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_1_Right_675
timestamp 1694700623
transform -1 0 17920 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_2_Left_513
timestamp 1694700623
transform 1 0 188272 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_2_Right_154
timestamp 1694700623
transform -1 0 204736 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_1_Left_335
timestamp 1694700623
transform 1 0 1344 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_1_Right_676
timestamp 1694700623
transform -1 0 17920 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_2_Left_514
timestamp 1694700623
transform 1 0 188272 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_2_Right_155
timestamp 1694700623
transform -1 0 204736 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_1_Left_336
timestamp 1694700623
transform 1 0 1344 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_1_Right_677
timestamp 1694700623
transform -1 0 17920 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_2_Left_515
timestamp 1694700623
transform 1 0 188272 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_2_Right_156
timestamp 1694700623
transform -1 0 204736 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_1_Left_337
timestamp 1694700623
transform 1 0 1344 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_1_Right_678
timestamp 1694700623
transform -1 0 17920 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_2_Left_516
timestamp 1694700623
transform 1 0 188272 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_2_Right_157
timestamp 1694700623
transform -1 0 204736 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_1_Left_338
timestamp 1694700623
transform 1 0 1344 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_1_Right_679
timestamp 1694700623
transform -1 0 17920 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_2_Left_517
timestamp 1694700623
transform 1 0 188272 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_2_Right_158
timestamp 1694700623
transform -1 0 204736 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_1_Left_339
timestamp 1694700623
transform 1 0 1344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_1_Right_680
timestamp 1694700623
transform -1 0 17920 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_2_Left_518
timestamp 1694700623
transform 1 0 188272 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_144_2_Right_159
timestamp 1694700623
transform -1 0 204736 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_1_Left_340
timestamp 1694700623
transform 1 0 1344 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_1_Right_681
timestamp 1694700623
transform -1 0 17920 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_2_Left_519
timestamp 1694700623
transform 1 0 188272 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_145_2_Right_160
timestamp 1694700623
transform -1 0 204736 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_1_Left_341
timestamp 1694700623
transform 1 0 1344 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_1_Right_682
timestamp 1694700623
transform -1 0 17920 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_2_Left_520
timestamp 1694700623
transform 1 0 188272 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_146_2_Right_161
timestamp 1694700623
transform -1 0 204736 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_1_Left_342
timestamp 1694700623
transform 1 0 1344 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_1_Right_683
timestamp 1694700623
transform -1 0 17920 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_2_Left_521
timestamp 1694700623
transform 1 0 188272 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_147_2_Right_162
timestamp 1694700623
transform -1 0 204736 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_1_Left_343
timestamp 1694700623
transform 1 0 1344 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_1_Right_684
timestamp 1694700623
transform -1 0 17920 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_2_Left_522
timestamp 1694700623
transform 1 0 188272 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_148_2_Right_163
timestamp 1694700623
transform -1 0 204736 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_149_1_Left_344
timestamp 1694700623
transform 1 0 1344 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_149_1_Right_685
timestamp 1694700623
transform -1 0 17920 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_149_2_Left_523
timestamp 1694700623
transform 1 0 188272 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_149_2_Right_164
timestamp 1694700623
transform -1 0 204736 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_150_1_Left_345
timestamp 1694700623
transform 1 0 1344 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_150_1_Right_686
timestamp 1694700623
transform -1 0 17920 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_150_2_Left_524
timestamp 1694700623
transform 1 0 188272 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_150_2_Right_165
timestamp 1694700623
transform -1 0 204736 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_151_1_Left_346
timestamp 1694700623
transform 1 0 1344 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_151_1_Right_687
timestamp 1694700623
transform -1 0 17920 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_151_2_Left_525
timestamp 1694700623
transform 1 0 188272 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_151_2_Right_166
timestamp 1694700623
transform -1 0 204736 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_152_1_Left_347
timestamp 1694700623
transform 1 0 1344 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_152_1_Right_688
timestamp 1694700623
transform -1 0 17920 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_152_2_Left_526
timestamp 1694700623
transform 1 0 188272 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_152_2_Right_167
timestamp 1694700623
transform -1 0 204736 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_153_1_Left_348
timestamp 1694700623
transform 1 0 1344 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_153_1_Right_689
timestamp 1694700623
transform -1 0 17920 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_153_2_Left_527
timestamp 1694700623
transform 1 0 188272 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_153_2_Right_168
timestamp 1694700623
transform -1 0 204736 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_154_1_Left_349
timestamp 1694700623
transform 1 0 1344 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_154_1_Right_690
timestamp 1694700623
transform -1 0 17920 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_154_2_Left_528
timestamp 1694700623
transform 1 0 188272 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_154_2_Right_169
timestamp 1694700623
transform -1 0 204736 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_155_1_Left_350
timestamp 1694700623
transform 1 0 1344 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_155_1_Right_691
timestamp 1694700623
transform -1 0 17920 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_155_2_Left_529
timestamp 1694700623
transform 1 0 188272 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_155_2_Right_170
timestamp 1694700623
transform -1 0 204736 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_156_1_Left_351
timestamp 1694700623
transform 1 0 1344 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_156_1_Right_692
timestamp 1694700623
transform -1 0 17920 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_156_2_Left_530
timestamp 1694700623
transform 1 0 188272 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_156_2_Right_171
timestamp 1694700623
transform -1 0 204736 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_157_1_Left_352
timestamp 1694700623
transform 1 0 1344 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_157_1_Right_693
timestamp 1694700623
transform -1 0 17920 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_157_2_Left_531
timestamp 1694700623
transform 1 0 188272 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_157_2_Right_172
timestamp 1694700623
transform -1 0 204736 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_158_1_Left_353
timestamp 1694700623
transform 1 0 1344 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_158_1_Right_694
timestamp 1694700623
transform -1 0 17920 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_158_2_Left_532
timestamp 1694700623
transform 1 0 188272 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_158_2_Right_173
timestamp 1694700623
transform -1 0 204736 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_159_1_Left_354
timestamp 1694700623
transform 1 0 1344 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_159_1_Right_695
timestamp 1694700623
transform -1 0 17920 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_159_2_Left_533
timestamp 1694700623
transform 1 0 188272 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_159_2_Right_174
timestamp 1694700623
transform -1 0 204736 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_160_1_Left_355
timestamp 1694700623
transform 1 0 1344 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_160_1_Right_696
timestamp 1694700623
transform -1 0 17920 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_160_2_Left_534
timestamp 1694700623
transform 1 0 188272 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_160_2_Right_175
timestamp 1694700623
transform -1 0 204736 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_161_1_Left_356
timestamp 1694700623
transform 1 0 1344 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_161_1_Right_697
timestamp 1694700623
transform -1 0 17920 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_161_2_Left_535
timestamp 1694700623
transform 1 0 188272 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_161_2_Right_176
timestamp 1694700623
transform -1 0 204736 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_162_1_Left_357
timestamp 1694700623
transform 1 0 1344 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_162_1_Right_698
timestamp 1694700623
transform -1 0 17920 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_162_2_Left_536
timestamp 1694700623
transform 1 0 188272 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_162_2_Right_177
timestamp 1694700623
transform -1 0 204736 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_163_1_Left_358
timestamp 1694700623
transform 1 0 1344 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_163_1_Right_699
timestamp 1694700623
transform -1 0 17920 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_163_2_Left_537
timestamp 1694700623
transform 1 0 188272 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_163_2_Right_178
timestamp 1694700623
transform -1 0 204736 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_164_1_Left_359
timestamp 1694700623
transform 1 0 1344 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_164_1_Right_700
timestamp 1694700623
transform -1 0 17920 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_164_2_Left_538
timestamp 1694700623
transform 1 0 188272 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_164_2_Right_179
timestamp 1694700623
transform -1 0 204736 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_165_1_Left_360
timestamp 1694700623
transform 1 0 1344 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_165_1_Right_701
timestamp 1694700623
transform -1 0 17920 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_165_2_Left_539
timestamp 1694700623
transform 1 0 188272 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_165_2_Right_180
timestamp 1694700623
transform -1 0 204736 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_166_1_Left_361
timestamp 1694700623
transform 1 0 1344 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_166_1_Right_702
timestamp 1694700623
transform -1 0 17920 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_166_2_Left_540
timestamp 1694700623
transform 1 0 188272 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_166_2_Right_181
timestamp 1694700623
transform -1 0 204736 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_167_1_Left_362
timestamp 1694700623
transform 1 0 1344 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_167_1_Right_703
timestamp 1694700623
transform -1 0 17920 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_167_2_Left_541
timestamp 1694700623
transform 1 0 188272 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_167_2_Right_182
timestamp 1694700623
transform -1 0 204736 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_168_1_Left_363
timestamp 1694700623
transform 1 0 1344 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_168_1_Right_704
timestamp 1694700623
transform -1 0 17920 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_168_2_Left_542
timestamp 1694700623
transform 1 0 188272 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_168_2_Right_183
timestamp 1694700623
transform -1 0 204736 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_169_1_Left_364
timestamp 1694700623
transform 1 0 1344 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_169_1_Right_705
timestamp 1694700623
transform -1 0 17920 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_169_2_Left_543
timestamp 1694700623
transform 1 0 188272 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_169_2_Right_184
timestamp 1694700623
transform -1 0 204736 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_170_1_Left_365
timestamp 1694700623
transform 1 0 1344 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_170_1_Right_706
timestamp 1694700623
transform -1 0 17920 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_170_2_Left_544
timestamp 1694700623
transform 1 0 188272 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_170_2_Right_185
timestamp 1694700623
transform -1 0 204736 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_171_1_Left_366
timestamp 1694700623
transform 1 0 1344 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_171_1_Right_707
timestamp 1694700623
transform -1 0 17920 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_171_2_Left_545
timestamp 1694700623
transform 1 0 188272 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_171_2_Right_186
timestamp 1694700623
transform -1 0 204736 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_172_1_Left_367
timestamp 1694700623
transform 1 0 1344 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_172_1_Right_708
timestamp 1694700623
transform -1 0 17920 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_172_2_Left_546
timestamp 1694700623
transform 1 0 188272 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_172_2_Right_187
timestamp 1694700623
transform -1 0 204736 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_173_1_Left_368
timestamp 1694700623
transform 1 0 1344 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_173_1_Right_709
timestamp 1694700623
transform -1 0 17920 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_173_2_Left_547
timestamp 1694700623
transform 1 0 188272 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_173_2_Right_188
timestamp 1694700623
transform -1 0 204736 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_174_1_Left_369
timestamp 1694700623
transform 1 0 1344 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_174_1_Right_710
timestamp 1694700623
transform -1 0 17920 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_174_2_Left_548
timestamp 1694700623
transform 1 0 188272 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_174_2_Right_189
timestamp 1694700623
transform -1 0 204736 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_175_1_Left_370
timestamp 1694700623
transform 1 0 1344 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_175_1_Right_711
timestamp 1694700623
transform -1 0 17920 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_175_2_Left_549
timestamp 1694700623
transform 1 0 188272 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_175_2_Right_190
timestamp 1694700623
transform -1 0 204736 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_176_1_Left_371
timestamp 1694700623
transform 1 0 1344 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_176_1_Right_712
timestamp 1694700623
transform -1 0 17920 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_176_2_Left_550
timestamp 1694700623
transform 1 0 188272 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_176_2_Right_191
timestamp 1694700623
transform -1 0 204736 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_177_1_Left_372
timestamp 1694700623
transform 1 0 1344 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_177_1_Right_713
timestamp 1694700623
transform -1 0 17920 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_177_2_Left_551
timestamp 1694700623
transform 1 0 188272 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_177_2_Right_192
timestamp 1694700623
transform -1 0 204736 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_178_1_Left_373
timestamp 1694700623
transform 1 0 1344 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_178_1_Right_714
timestamp 1694700623
transform -1 0 17920 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_178_2_Left_552
timestamp 1694700623
transform 1 0 188272 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_178_2_Right_193
timestamp 1694700623
transform -1 0 204736 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_179_1_Left_374
timestamp 1694700623
transform 1 0 1344 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_179_1_Right_715
timestamp 1694700623
transform -1 0 17920 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_179_2_Left_553
timestamp 1694700623
transform 1 0 188272 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_179_2_Right_194
timestamp 1694700623
transform -1 0 204736 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_180_1_Left_375
timestamp 1694700623
transform 1 0 1344 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_180_1_Right_716
timestamp 1694700623
transform -1 0 17920 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_180_2_Left_554
timestamp 1694700623
transform 1 0 188272 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_180_2_Right_195
timestamp 1694700623
transform -1 0 204736 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_181_Left_376
timestamp 1694700623
transform 1 0 1344 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_181_Right_18
timestamp 1694700623
transform -1 0 204736 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_182_Left_377
timestamp 1694700623
transform 1 0 1344 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_182_Right_19
timestamp 1694700623
transform -1 0 204736 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_183_Left_378
timestamp 1694700623
transform 1 0 1344 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_183_Right_20
timestamp 1694700623
transform -1 0 204736 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_184_Left_379
timestamp 1694700623
transform 1 0 1344 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_184_Right_21
timestamp 1694700623
transform -1 0 204736 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_185_Left_380
timestamp 1694700623
transform 1 0 1344 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_185_Right_22
timestamp 1694700623
transform -1 0 204736 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_186_Left_381
timestamp 1694700623
transform 1 0 1344 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_186_Right_23
timestamp 1694700623
transform -1 0 204736 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_187_Left_382
timestamp 1694700623
transform 1 0 1344 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_187_Right_24
timestamp 1694700623
transform -1 0 204736 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_188_Left_383
timestamp 1694700623
transform 1 0 1344 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_188_Right_25
timestamp 1694700623
transform -1 0 204736 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_189_Left_384
timestamp 1694700623
transform 1 0 1344 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_189_Right_26
timestamp 1694700623
transform -1 0 204736 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_190_Left_385
timestamp 1694700623
transform 1 0 1344 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_190_Right_27
timestamp 1694700623
transform -1 0 204736 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_191_Left_386
timestamp 1694700623
transform 1 0 1344 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_191_Right_28
timestamp 1694700623
transform -1 0 204736 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_192_Left_387
timestamp 1694700623
transform 1 0 1344 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_192_Right_29
timestamp 1694700623
transform -1 0 204736 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_193_Left_388
timestamp 1694700623
transform 1 0 1344 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_193_Right_30
timestamp 1694700623
transform -1 0 204736 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_194_Left_389
timestamp 1694700623
transform 1 0 1344 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_194_Right_31
timestamp 1694700623
transform -1 0 204736 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_195_Left_390
timestamp 1694700623
transform 1 0 1344 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_195_Right_32
timestamp 1694700623
transform -1 0 204736 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_718 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_719
timestamp 1694700623
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_720
timestamp 1694700623
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_721
timestamp 1694700623
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_722
timestamp 1694700623
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_723
timestamp 1694700623
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_724
timestamp 1694700623
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_725
timestamp 1694700623
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_726
timestamp 1694700623
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_727
timestamp 1694700623
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_728
timestamp 1694700623
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_729
timestamp 1694700623
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_730
timestamp 1694700623
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_731
timestamp 1694700623
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_732
timestamp 1694700623
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_733
timestamp 1694700623
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_734
timestamp 1694700623
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_735
timestamp 1694700623
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_736
timestamp 1694700623
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_737
timestamp 1694700623
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_738
timestamp 1694700623
transform 1 0 81312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_739
timestamp 1694700623
transform 1 0 85120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_740
timestamp 1694700623
transform 1 0 88928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_741
timestamp 1694700623
transform 1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_742
timestamp 1694700623
transform 1 0 96544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_743
timestamp 1694700623
transform 1 0 100352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_744
timestamp 1694700623
transform 1 0 104160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_745
timestamp 1694700623
transform 1 0 107968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_746
timestamp 1694700623
transform 1 0 111776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_747
timestamp 1694700623
transform 1 0 115584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_748
timestamp 1694700623
transform 1 0 119392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_749
timestamp 1694700623
transform 1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_750
timestamp 1694700623
transform 1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_751
timestamp 1694700623
transform 1 0 130816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_752
timestamp 1694700623
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_753
timestamp 1694700623
transform 1 0 138432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_754
timestamp 1694700623
transform 1 0 142240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_755
timestamp 1694700623
transform 1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_756
timestamp 1694700623
transform 1 0 149856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_757
timestamp 1694700623
transform 1 0 153664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_758
timestamp 1694700623
transform 1 0 157472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_759
timestamp 1694700623
transform 1 0 161280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_760
timestamp 1694700623
transform 1 0 165088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_761
timestamp 1694700623
transform 1 0 168896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_762
timestamp 1694700623
transform 1 0 172704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_763
timestamp 1694700623
transform 1 0 176512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_764
timestamp 1694700623
transform 1 0 180320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_765
timestamp 1694700623
transform 1 0 184128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_766
timestamp 1694700623
transform 1 0 187936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_767
timestamp 1694700623
transform 1 0 191744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_768
timestamp 1694700623
transform 1 0 195552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_769
timestamp 1694700623
transform 1 0 199360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_770
timestamp 1694700623
transform 1 0 203168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_771
timestamp 1694700623
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_772
timestamp 1694700623
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_773
timestamp 1694700623
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_774
timestamp 1694700623
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_775
timestamp 1694700623
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_776
timestamp 1694700623
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_777
timestamp 1694700623
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_778
timestamp 1694700623
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_779
timestamp 1694700623
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_780
timestamp 1694700623
transform 1 0 79744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_781
timestamp 1694700623
transform 1 0 87584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_782
timestamp 1694700623
transform 1 0 95424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_783
timestamp 1694700623
transform 1 0 103264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_784
timestamp 1694700623
transform 1 0 111104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_785
timestamp 1694700623
transform 1 0 118944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_786
timestamp 1694700623
transform 1 0 126784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_787
timestamp 1694700623
transform 1 0 134624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_788
timestamp 1694700623
transform 1 0 142464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_789
timestamp 1694700623
transform 1 0 150304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_790
timestamp 1694700623
transform 1 0 158144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_791
timestamp 1694700623
transform 1 0 165984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_792
timestamp 1694700623
transform 1 0 173824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_793
timestamp 1694700623
transform 1 0 181664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_794
timestamp 1694700623
transform 1 0 189504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_795
timestamp 1694700623
transform 1 0 197344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_796
timestamp 1694700623
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_797
timestamp 1694700623
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_798
timestamp 1694700623
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_799
timestamp 1694700623
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_800
timestamp 1694700623
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_801
timestamp 1694700623
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_802
timestamp 1694700623
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_803
timestamp 1694700623
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_804
timestamp 1694700623
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_805
timestamp 1694700623
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_806
timestamp 1694700623
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_807
timestamp 1694700623
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_808
timestamp 1694700623
transform 1 0 99344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_809
timestamp 1694700623
transform 1 0 107184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_810
timestamp 1694700623
transform 1 0 115024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_811
timestamp 1694700623
transform 1 0 122864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_812
timestamp 1694700623
transform 1 0 130704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_813
timestamp 1694700623
transform 1 0 138544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_814
timestamp 1694700623
transform 1 0 146384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_815
timestamp 1694700623
transform 1 0 154224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_816
timestamp 1694700623
transform 1 0 162064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_817
timestamp 1694700623
transform 1 0 169904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_818
timestamp 1694700623
transform 1 0 177744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_819
timestamp 1694700623
transform 1 0 185584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_820
timestamp 1694700623
transform 1 0 193424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_821
timestamp 1694700623
transform 1 0 201264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_822
timestamp 1694700623
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_823
timestamp 1694700623
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_824
timestamp 1694700623
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_825
timestamp 1694700623
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_826
timestamp 1694700623
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_827
timestamp 1694700623
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_828
timestamp 1694700623
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_829
timestamp 1694700623
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_830
timestamp 1694700623
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_831
timestamp 1694700623
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_832
timestamp 1694700623
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_833
timestamp 1694700623
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_834
timestamp 1694700623
transform 1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_835
timestamp 1694700623
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_836
timestamp 1694700623
transform 1 0 118944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_837
timestamp 1694700623
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_838
timestamp 1694700623
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_839
timestamp 1694700623
transform 1 0 142464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_840
timestamp 1694700623
transform 1 0 150304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_841
timestamp 1694700623
transform 1 0 158144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_842
timestamp 1694700623
transform 1 0 165984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_843
timestamp 1694700623
transform 1 0 173824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_844
timestamp 1694700623
transform 1 0 181664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_845
timestamp 1694700623
transform 1 0 189504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_846
timestamp 1694700623
transform 1 0 197344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_847
timestamp 1694700623
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_848
timestamp 1694700623
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_849
timestamp 1694700623
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_850
timestamp 1694700623
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_851
timestamp 1694700623
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_852
timestamp 1694700623
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_853
timestamp 1694700623
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_854
timestamp 1694700623
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_855
timestamp 1694700623
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_856
timestamp 1694700623
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_857
timestamp 1694700623
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_858
timestamp 1694700623
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_859
timestamp 1694700623
transform 1 0 99344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_860
timestamp 1694700623
transform 1 0 107184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_861
timestamp 1694700623
transform 1 0 115024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_862
timestamp 1694700623
transform 1 0 122864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_863
timestamp 1694700623
transform 1 0 130704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_864
timestamp 1694700623
transform 1 0 138544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_865
timestamp 1694700623
transform 1 0 146384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_866
timestamp 1694700623
transform 1 0 154224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_867
timestamp 1694700623
transform 1 0 162064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_868
timestamp 1694700623
transform 1 0 169904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_869
timestamp 1694700623
transform 1 0 177744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_870
timestamp 1694700623
transform 1 0 185584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_871
timestamp 1694700623
transform 1 0 193424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_872
timestamp 1694700623
transform 1 0 201264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_873
timestamp 1694700623
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_874
timestamp 1694700623
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_875
timestamp 1694700623
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_876
timestamp 1694700623
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_877
timestamp 1694700623
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_878
timestamp 1694700623
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_879
timestamp 1694700623
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_880
timestamp 1694700623
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_881
timestamp 1694700623
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_882
timestamp 1694700623
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_883
timestamp 1694700623
transform 1 0 87584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_884
timestamp 1694700623
transform 1 0 95424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_885
timestamp 1694700623
transform 1 0 103264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_886
timestamp 1694700623
transform 1 0 111104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_887
timestamp 1694700623
transform 1 0 118944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_888
timestamp 1694700623
transform 1 0 126784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_889
timestamp 1694700623
transform 1 0 134624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_890
timestamp 1694700623
transform 1 0 142464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_891
timestamp 1694700623
transform 1 0 150304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_892
timestamp 1694700623
transform 1 0 158144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_893
timestamp 1694700623
transform 1 0 165984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_894
timestamp 1694700623
transform 1 0 173824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_895
timestamp 1694700623
transform 1 0 181664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_896
timestamp 1694700623
transform 1 0 189504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_897
timestamp 1694700623
transform 1 0 197344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_898
timestamp 1694700623
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_899
timestamp 1694700623
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_900
timestamp 1694700623
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_901
timestamp 1694700623
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_902
timestamp 1694700623
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_903
timestamp 1694700623
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_904
timestamp 1694700623
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_905
timestamp 1694700623
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_906
timestamp 1694700623
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_907
timestamp 1694700623
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_908
timestamp 1694700623
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_909
timestamp 1694700623
transform 1 0 91504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_910
timestamp 1694700623
transform 1 0 99344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_911
timestamp 1694700623
transform 1 0 107184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_912
timestamp 1694700623
transform 1 0 115024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_913
timestamp 1694700623
transform 1 0 122864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_914
timestamp 1694700623
transform 1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_915
timestamp 1694700623
transform 1 0 138544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_916
timestamp 1694700623
transform 1 0 146384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_917
timestamp 1694700623
transform 1 0 154224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_918
timestamp 1694700623
transform 1 0 162064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_919
timestamp 1694700623
transform 1 0 169904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_920
timestamp 1694700623
transform 1 0 177744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_921
timestamp 1694700623
transform 1 0 185584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_922
timestamp 1694700623
transform 1 0 193424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_923
timestamp 1694700623
transform 1 0 201264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_924
timestamp 1694700623
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_925
timestamp 1694700623
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_926
timestamp 1694700623
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_927
timestamp 1694700623
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_928
timestamp 1694700623
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_929
timestamp 1694700623
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_930
timestamp 1694700623
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_931
timestamp 1694700623
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_932
timestamp 1694700623
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_933
timestamp 1694700623
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_934
timestamp 1694700623
transform 1 0 87584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_935
timestamp 1694700623
transform 1 0 95424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_936
timestamp 1694700623
transform 1 0 103264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_937
timestamp 1694700623
transform 1 0 111104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_938
timestamp 1694700623
transform 1 0 118944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_939
timestamp 1694700623
transform 1 0 126784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_940
timestamp 1694700623
transform 1 0 134624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_941
timestamp 1694700623
transform 1 0 142464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_942
timestamp 1694700623
transform 1 0 150304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_943
timestamp 1694700623
transform 1 0 158144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_944
timestamp 1694700623
transform 1 0 165984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_945
timestamp 1694700623
transform 1 0 173824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_946
timestamp 1694700623
transform 1 0 181664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_947
timestamp 1694700623
transform 1 0 189504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_948
timestamp 1694700623
transform 1 0 197344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_949
timestamp 1694700623
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_950
timestamp 1694700623
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_951
timestamp 1694700623
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_952
timestamp 1694700623
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_953
timestamp 1694700623
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_954
timestamp 1694700623
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_955
timestamp 1694700623
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_956
timestamp 1694700623
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_957
timestamp 1694700623
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_958
timestamp 1694700623
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_959
timestamp 1694700623
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_960
timestamp 1694700623
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_961
timestamp 1694700623
transform 1 0 99344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_962
timestamp 1694700623
transform 1 0 107184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_963
timestamp 1694700623
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_964
timestamp 1694700623
transform 1 0 122864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_965
timestamp 1694700623
transform 1 0 130704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_966
timestamp 1694700623
transform 1 0 138544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_967
timestamp 1694700623
transform 1 0 146384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_968
timestamp 1694700623
transform 1 0 154224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_969
timestamp 1694700623
transform 1 0 162064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_970
timestamp 1694700623
transform 1 0 169904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_971
timestamp 1694700623
transform 1 0 177744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_972
timestamp 1694700623
transform 1 0 185584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_973
timestamp 1694700623
transform 1 0 193424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_974
timestamp 1694700623
transform 1 0 201264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_975
timestamp 1694700623
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_976
timestamp 1694700623
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_977
timestamp 1694700623
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_978
timestamp 1694700623
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_979
timestamp 1694700623
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_980
timestamp 1694700623
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_981
timestamp 1694700623
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_982
timestamp 1694700623
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_983
timestamp 1694700623
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_984
timestamp 1694700623
transform 1 0 79744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_985
timestamp 1694700623
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_986
timestamp 1694700623
transform 1 0 95424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_987
timestamp 1694700623
transform 1 0 103264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_988
timestamp 1694700623
transform 1 0 111104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_989
timestamp 1694700623
transform 1 0 118944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_990
timestamp 1694700623
transform 1 0 126784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_991
timestamp 1694700623
transform 1 0 134624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_992
timestamp 1694700623
transform 1 0 142464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_993
timestamp 1694700623
transform 1 0 150304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_994
timestamp 1694700623
transform 1 0 158144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_995
timestamp 1694700623
transform 1 0 165984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_996
timestamp 1694700623
transform 1 0 173824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_997
timestamp 1694700623
transform 1 0 181664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_998
timestamp 1694700623
transform 1 0 189504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_999
timestamp 1694700623
transform 1 0 197344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1000
timestamp 1694700623
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1001
timestamp 1694700623
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1002
timestamp 1694700623
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1003
timestamp 1694700623
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1004
timestamp 1694700623
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1005
timestamp 1694700623
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1006
timestamp 1694700623
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1007
timestamp 1694700623
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1008
timestamp 1694700623
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1009
timestamp 1694700623
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1010
timestamp 1694700623
transform 1 0 83664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1011
timestamp 1694700623
transform 1 0 91504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1012
timestamp 1694700623
transform 1 0 99344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1013
timestamp 1694700623
transform 1 0 107184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1014
timestamp 1694700623
transform 1 0 115024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1015
timestamp 1694700623
transform 1 0 122864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1016
timestamp 1694700623
transform 1 0 130704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1017
timestamp 1694700623
transform 1 0 138544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1018
timestamp 1694700623
transform 1 0 146384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1019
timestamp 1694700623
transform 1 0 154224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1020
timestamp 1694700623
transform 1 0 162064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1021
timestamp 1694700623
transform 1 0 169904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1022
timestamp 1694700623
transform 1 0 177744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1023
timestamp 1694700623
transform 1 0 185584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1024
timestamp 1694700623
transform 1 0 193424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_1025
timestamp 1694700623
transform 1 0 201264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1026
timestamp 1694700623
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1027
timestamp 1694700623
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1028
timestamp 1694700623
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1029
timestamp 1694700623
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1030
timestamp 1694700623
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1031
timestamp 1694700623
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1032
timestamp 1694700623
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1033
timestamp 1694700623
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1034
timestamp 1694700623
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1035
timestamp 1694700623
transform 1 0 79744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1036
timestamp 1694700623
transform 1 0 87584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1037
timestamp 1694700623
transform 1 0 95424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1038
timestamp 1694700623
transform 1 0 103264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1039
timestamp 1694700623
transform 1 0 111104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1040
timestamp 1694700623
transform 1 0 118944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1041
timestamp 1694700623
transform 1 0 126784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1042
timestamp 1694700623
transform 1 0 134624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1043
timestamp 1694700623
transform 1 0 142464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1044
timestamp 1694700623
transform 1 0 150304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1045
timestamp 1694700623
transform 1 0 158144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1046
timestamp 1694700623
transform 1 0 165984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1047
timestamp 1694700623
transform 1 0 173824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1048
timestamp 1694700623
transform 1 0 181664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1049
timestamp 1694700623
transform 1 0 189504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_1050
timestamp 1694700623
transform 1 0 197344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1051
timestamp 1694700623
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1052
timestamp 1694700623
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1053
timestamp 1694700623
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1054
timestamp 1694700623
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1055
timestamp 1694700623
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1056
timestamp 1694700623
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1057
timestamp 1694700623
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1058
timestamp 1694700623
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1059
timestamp 1694700623
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1060
timestamp 1694700623
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1061
timestamp 1694700623
transform 1 0 83664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1062
timestamp 1694700623
transform 1 0 91504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1063
timestamp 1694700623
transform 1 0 99344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1064
timestamp 1694700623
transform 1 0 107184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1065
timestamp 1694700623
transform 1 0 115024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1066
timestamp 1694700623
transform 1 0 122864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1067
timestamp 1694700623
transform 1 0 130704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1068
timestamp 1694700623
transform 1 0 138544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1069
timestamp 1694700623
transform 1 0 146384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1070
timestamp 1694700623
transform 1 0 154224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1071
timestamp 1694700623
transform 1 0 162064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1072
timestamp 1694700623
transform 1 0 169904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1073
timestamp 1694700623
transform 1 0 177744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1074
timestamp 1694700623
transform 1 0 185584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1075
timestamp 1694700623
transform 1 0 193424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_1076
timestamp 1694700623
transform 1 0 201264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1077
timestamp 1694700623
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1078
timestamp 1694700623
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1079
timestamp 1694700623
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1080
timestamp 1694700623
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1081
timestamp 1694700623
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1082
timestamp 1694700623
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1083
timestamp 1694700623
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1084
timestamp 1694700623
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1085
timestamp 1694700623
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1086
timestamp 1694700623
transform 1 0 79744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1087
timestamp 1694700623
transform 1 0 87584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1088
timestamp 1694700623
transform 1 0 95424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1089
timestamp 1694700623
transform 1 0 103264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1090
timestamp 1694700623
transform 1 0 111104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1091
timestamp 1694700623
transform 1 0 118944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1092
timestamp 1694700623
transform 1 0 126784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1093
timestamp 1694700623
transform 1 0 134624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1094
timestamp 1694700623
transform 1 0 142464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1095
timestamp 1694700623
transform 1 0 150304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1096
timestamp 1694700623
transform 1 0 158144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1097
timestamp 1694700623
transform 1 0 165984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1098
timestamp 1694700623
transform 1 0 173824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1099
timestamp 1694700623
transform 1 0 181664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1100
timestamp 1694700623
transform 1 0 189504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_1101
timestamp 1694700623
transform 1 0 197344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1102
timestamp 1694700623
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1103
timestamp 1694700623
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1104
timestamp 1694700623
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1105
timestamp 1694700623
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1106
timestamp 1694700623
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1107
timestamp 1694700623
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1108
timestamp 1694700623
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1109
timestamp 1694700623
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1110
timestamp 1694700623
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1111
timestamp 1694700623
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1112
timestamp 1694700623
transform 1 0 83664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1113
timestamp 1694700623
transform 1 0 91504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1114
timestamp 1694700623
transform 1 0 99344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1115
timestamp 1694700623
transform 1 0 107184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1116
timestamp 1694700623
transform 1 0 115024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1117
timestamp 1694700623
transform 1 0 122864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1118
timestamp 1694700623
transform 1 0 130704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1119
timestamp 1694700623
transform 1 0 138544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1120
timestamp 1694700623
transform 1 0 146384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1121
timestamp 1694700623
transform 1 0 154224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1122
timestamp 1694700623
transform 1 0 162064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1123
timestamp 1694700623
transform 1 0 169904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1124
timestamp 1694700623
transform 1 0 177744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1125
timestamp 1694700623
transform 1 0 185584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1126
timestamp 1694700623
transform 1 0 193424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_1127
timestamp 1694700623
transform 1 0 201264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1128
timestamp 1694700623
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1129
timestamp 1694700623
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1130
timestamp 1694700623
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1131
timestamp 1694700623
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1132
timestamp 1694700623
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1133
timestamp 1694700623
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1134
timestamp 1694700623
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1135
timestamp 1694700623
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1136
timestamp 1694700623
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1137
timestamp 1694700623
transform 1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1138
timestamp 1694700623
transform 1 0 87584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1139
timestamp 1694700623
transform 1 0 95424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1140
timestamp 1694700623
transform 1 0 103264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1141
timestamp 1694700623
transform 1 0 111104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1142
timestamp 1694700623
transform 1 0 118944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1143
timestamp 1694700623
transform 1 0 126784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1144
timestamp 1694700623
transform 1 0 134624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1145
timestamp 1694700623
transform 1 0 142464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1146
timestamp 1694700623
transform 1 0 150304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1147
timestamp 1694700623
transform 1 0 158144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1148
timestamp 1694700623
transform 1 0 165984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1149
timestamp 1694700623
transform 1 0 173824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1150
timestamp 1694700623
transform 1 0 181664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1151
timestamp 1694700623
transform 1 0 189504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_1152
timestamp 1694700623
transform 1 0 197344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1153
timestamp 1694700623
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1154
timestamp 1694700623
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1155
timestamp 1694700623
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1156
timestamp 1694700623
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1157
timestamp 1694700623
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1158
timestamp 1694700623
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1159
timestamp 1694700623
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1160
timestamp 1694700623
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1161
timestamp 1694700623
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1162
timestamp 1694700623
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1163
timestamp 1694700623
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1164
timestamp 1694700623
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1165
timestamp 1694700623
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1166
timestamp 1694700623
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1167
timestamp 1694700623
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1168
timestamp 1694700623
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1169
timestamp 1694700623
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1170
timestamp 1694700623
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1171
timestamp 1694700623
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1172
timestamp 1694700623
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1173
timestamp 1694700623
transform 1 0 162064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1174
timestamp 1694700623
transform 1 0 169904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1175
timestamp 1694700623
transform 1 0 177744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1176
timestamp 1694700623
transform 1 0 185584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1177
timestamp 1694700623
transform 1 0 193424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_1178
timestamp 1694700623
transform 1 0 201264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1179
timestamp 1694700623
transform 1 0 5152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1180
timestamp 1694700623
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1181
timestamp 1694700623
transform 1 0 12768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1182
timestamp 1694700623
transform 1 0 16576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1183
timestamp 1694700623
transform 1 0 20384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1184
timestamp 1694700623
transform 1 0 24192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1185
timestamp 1694700623
transform 1 0 28000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1186
timestamp 1694700623
transform 1 0 31808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1187
timestamp 1694700623
transform 1 0 35616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1188
timestamp 1694700623
transform 1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1189
timestamp 1694700623
transform 1 0 43232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1190
timestamp 1694700623
transform 1 0 47040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1191
timestamp 1694700623
transform 1 0 50848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1192
timestamp 1694700623
transform 1 0 54656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1193
timestamp 1694700623
transform 1 0 58464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1194
timestamp 1694700623
transform 1 0 62272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1195
timestamp 1694700623
transform 1 0 66080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1196
timestamp 1694700623
transform 1 0 69888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1197
timestamp 1694700623
transform 1 0 73696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1198
timestamp 1694700623
transform 1 0 77504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1199
timestamp 1694700623
transform 1 0 81312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1200
timestamp 1694700623
transform 1 0 85120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1201
timestamp 1694700623
transform 1 0 88928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1202
timestamp 1694700623
transform 1 0 92736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1203
timestamp 1694700623
transform 1 0 96544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1204
timestamp 1694700623
transform 1 0 100352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1205
timestamp 1694700623
transform 1 0 104160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1206
timestamp 1694700623
transform 1 0 107968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1207
timestamp 1694700623
transform 1 0 111776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1208
timestamp 1694700623
transform 1 0 115584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1209
timestamp 1694700623
transform 1 0 119392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1210
timestamp 1694700623
transform 1 0 123200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1211
timestamp 1694700623
transform 1 0 127008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1212
timestamp 1694700623
transform 1 0 130816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1213
timestamp 1694700623
transform 1 0 134624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1214
timestamp 1694700623
transform 1 0 138432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1215
timestamp 1694700623
transform 1 0 142240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1216
timestamp 1694700623
transform 1 0 146048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1217
timestamp 1694700623
transform 1 0 149856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1218
timestamp 1694700623
transform 1 0 153664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1219
timestamp 1694700623
transform 1 0 157472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1220
timestamp 1694700623
transform 1 0 161280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1221
timestamp 1694700623
transform 1 0 165088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1222
timestamp 1694700623
transform 1 0 168896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1223
timestamp 1694700623
transform 1 0 172704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1224
timestamp 1694700623
transform 1 0 176512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1225
timestamp 1694700623
transform 1 0 180320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1226
timestamp 1694700623
transform 1 0 184128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1227
timestamp 1694700623
transform 1 0 187936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1228
timestamp 1694700623
transform 1 0 191744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1229
timestamp 1694700623
transform 1 0 195552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1230
timestamp 1694700623
transform 1 0 199360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_1231
timestamp 1694700623
transform 1 0 203168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_1_1994
timestamp 1694700623
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_1_1995
timestamp 1694700623
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_2_1996
timestamp 1694700623
transform 1 0 192192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_2_1997
timestamp 1694700623
transform 1 0 200032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_1_1232
timestamp 1694700623
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_1_1233
timestamp 1694700623
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_2_1998
timestamp 1694700623
transform 1 0 196112 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_2_1999
timestamp 1694700623
transform 1 0 203952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_1_1234
timestamp 1694700623
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_1_1235
timestamp 1694700623
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_2_2000
timestamp 1694700623
transform 1 0 192192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_2_2001
timestamp 1694700623
transform 1 0 200032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_1_1236
timestamp 1694700623
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_1_1237
timestamp 1694700623
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_2_2002
timestamp 1694700623
transform 1 0 196112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_2_2003
timestamp 1694700623
transform 1 0 203952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1_1238
timestamp 1694700623
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_1_1239
timestamp 1694700623
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_2_2004
timestamp 1694700623
transform 1 0 192192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_2_2005
timestamp 1694700623
transform 1 0 200032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1_1240
timestamp 1694700623
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_1_1241
timestamp 1694700623
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_2_2006
timestamp 1694700623
transform 1 0 196112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_2_2007
timestamp 1694700623
transform 1 0 203952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1_1242
timestamp 1694700623
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_1_1243
timestamp 1694700623
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_2_2008
timestamp 1694700623
transform 1 0 192192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_2_2009
timestamp 1694700623
transform 1 0 200032 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1_1244
timestamp 1694700623
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_1_1245
timestamp 1694700623
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_2_2010
timestamp 1694700623
transform 1 0 196112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_2_2011
timestamp 1694700623
transform 1 0 203952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1_1246
timestamp 1694700623
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_1_1247
timestamp 1694700623
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_2_2012
timestamp 1694700623
transform 1 0 192192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_2_2013
timestamp 1694700623
transform 1 0 200032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1_1248
timestamp 1694700623
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_1_1249
timestamp 1694700623
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_2_2014
timestamp 1694700623
transform 1 0 196112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_2_2015
timestamp 1694700623
transform 1 0 203952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1_1250
timestamp 1694700623
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_1_1251
timestamp 1694700623
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_2_2016
timestamp 1694700623
transform 1 0 192192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_2_2017
timestamp 1694700623
transform 1 0 200032 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1_1252
timestamp 1694700623
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_1_1253
timestamp 1694700623
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_2_2018
timestamp 1694700623
transform 1 0 196112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_2_2019
timestamp 1694700623
transform 1 0 203952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1_1254
timestamp 1694700623
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_1_1255
timestamp 1694700623
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_2_2020
timestamp 1694700623
transform 1 0 192192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_2_2021
timestamp 1694700623
transform 1 0 200032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1_1256
timestamp 1694700623
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1_1257
timestamp 1694700623
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_2_2022
timestamp 1694700623
transform 1 0 196112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_2_2023
timestamp 1694700623
transform 1 0 203952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1_1258
timestamp 1694700623
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1_1259
timestamp 1694700623
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_2_2024
timestamp 1694700623
transform 1 0 192192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_2_2025
timestamp 1694700623
transform 1 0 200032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1_1260
timestamp 1694700623
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1_1261
timestamp 1694700623
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_2_2026
timestamp 1694700623
transform 1 0 196112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_2_2027
timestamp 1694700623
transform 1 0 203952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1_1262
timestamp 1694700623
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1_1263
timestamp 1694700623
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_2_2028
timestamp 1694700623
transform 1 0 192192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_2_2029
timestamp 1694700623
transform 1 0 200032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1_1264
timestamp 1694700623
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1_1265
timestamp 1694700623
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_2_2030
timestamp 1694700623
transform 1 0 196112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_2_2031
timestamp 1694700623
transform 1 0 203952 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1_1266
timestamp 1694700623
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1_1267
timestamp 1694700623
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_2_2032
timestamp 1694700623
transform 1 0 192192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_2_2033
timestamp 1694700623
transform 1 0 200032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1_1268
timestamp 1694700623
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1_1269
timestamp 1694700623
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_2_2034
timestamp 1694700623
transform 1 0 196112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_2_2035
timestamp 1694700623
transform 1 0 203952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1_1270
timestamp 1694700623
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1_1271
timestamp 1694700623
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_2_2036
timestamp 1694700623
transform 1 0 192192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_2_2037
timestamp 1694700623
transform 1 0 200032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1_1272
timestamp 1694700623
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1_1273
timestamp 1694700623
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_2_2038
timestamp 1694700623
transform 1 0 196112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_2_2039
timestamp 1694700623
transform 1 0 203952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1_1274
timestamp 1694700623
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1_1275
timestamp 1694700623
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_2_2040
timestamp 1694700623
transform 1 0 192192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_2_2041
timestamp 1694700623
transform 1 0 200032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1_1276
timestamp 1694700623
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1_1277
timestamp 1694700623
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_2_2042
timestamp 1694700623
transform 1 0 196112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_2_2043
timestamp 1694700623
transform 1 0 203952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1_1278
timestamp 1694700623
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1_1279
timestamp 1694700623
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_2_2044
timestamp 1694700623
transform 1 0 192192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_2_2045
timestamp 1694700623
transform 1 0 200032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1_1280
timestamp 1694700623
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1_1281
timestamp 1694700623
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_2_2046
timestamp 1694700623
transform 1 0 196112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_2_2047
timestamp 1694700623
transform 1 0 203952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1_1282
timestamp 1694700623
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1_1283
timestamp 1694700623
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_2_2048
timestamp 1694700623
transform 1 0 192192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_2_2049
timestamp 1694700623
transform 1 0 200032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1_1284
timestamp 1694700623
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1_1285
timestamp 1694700623
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_2_2050
timestamp 1694700623
transform 1 0 196112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_2_2051
timestamp 1694700623
transform 1 0 203952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1_1286
timestamp 1694700623
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1_1287
timestamp 1694700623
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_2_2052
timestamp 1694700623
transform 1 0 192192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_2_2053
timestamp 1694700623
transform 1 0 200032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1_1288
timestamp 1694700623
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1_1289
timestamp 1694700623
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_2_2054
timestamp 1694700623
transform 1 0 196112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_2_2055
timestamp 1694700623
transform 1 0 203952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1_1290
timestamp 1694700623
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1_1291
timestamp 1694700623
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2_2056
timestamp 1694700623
transform 1 0 192192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_2_2057
timestamp 1694700623
transform 1 0 200032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1_1292
timestamp 1694700623
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1_1293
timestamp 1694700623
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2_2058
timestamp 1694700623
transform 1 0 196112 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_2_2059
timestamp 1694700623
transform 1 0 203952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1_1294
timestamp 1694700623
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1_1295
timestamp 1694700623
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2_2060
timestamp 1694700623
transform 1 0 192192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_2_2061
timestamp 1694700623
transform 1 0 200032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1_1296
timestamp 1694700623
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1_1297
timestamp 1694700623
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2_2062
timestamp 1694700623
transform 1 0 196112 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_2_2063
timestamp 1694700623
transform 1 0 203952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1_1298
timestamp 1694700623
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1_1299
timestamp 1694700623
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2_2064
timestamp 1694700623
transform 1 0 192192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_2_2065
timestamp 1694700623
transform 1 0 200032 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1_1300
timestamp 1694700623
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1_1301
timestamp 1694700623
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2_2066
timestamp 1694700623
transform 1 0 196112 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_2_2067
timestamp 1694700623
transform 1 0 203952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1_1302
timestamp 1694700623
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1_1303
timestamp 1694700623
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2_2068
timestamp 1694700623
transform 1 0 192192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_2_2069
timestamp 1694700623
transform 1 0 200032 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1_1304
timestamp 1694700623
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_1_1305
timestamp 1694700623
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2_2070
timestamp 1694700623
transform 1 0 196112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_2_2071
timestamp 1694700623
transform 1 0 203952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1_1306
timestamp 1694700623
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_1_1307
timestamp 1694700623
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2_2072
timestamp 1694700623
transform 1 0 192192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_2_2073
timestamp 1694700623
transform 1 0 200032 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1_1308
timestamp 1694700623
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_1_1309
timestamp 1694700623
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2_2074
timestamp 1694700623
transform 1 0 196112 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_2_2075
timestamp 1694700623
transform 1 0 203952 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1_1310
timestamp 1694700623
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_1_1311
timestamp 1694700623
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2_2076
timestamp 1694700623
transform 1 0 192192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_2_2077
timestamp 1694700623
transform 1 0 200032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1_1312
timestamp 1694700623
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_1_1313
timestamp 1694700623
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2_2078
timestamp 1694700623
transform 1 0 196112 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_2_2079
timestamp 1694700623
transform 1 0 203952 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1_1314
timestamp 1694700623
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_1_1315
timestamp 1694700623
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2_2080
timestamp 1694700623
transform 1 0 192192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_2_2081
timestamp 1694700623
transform 1 0 200032 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1_1316
timestamp 1694700623
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_1_1317
timestamp 1694700623
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2_2082
timestamp 1694700623
transform 1 0 196112 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_2_2083
timestamp 1694700623
transform 1 0 203952 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1_1318
timestamp 1694700623
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_1_1319
timestamp 1694700623
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2_2084
timestamp 1694700623
transform 1 0 192192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_2_2085
timestamp 1694700623
transform 1 0 200032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1_1320
timestamp 1694700623
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_1_1321
timestamp 1694700623
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2_2086
timestamp 1694700623
transform 1 0 196112 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_2_2087
timestamp 1694700623
transform 1 0 203952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1_1322
timestamp 1694700623
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_1_1323
timestamp 1694700623
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2_2088
timestamp 1694700623
transform 1 0 192192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_2_2089
timestamp 1694700623
transform 1 0 200032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1_1324
timestamp 1694700623
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_1_1325
timestamp 1694700623
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2_2090
timestamp 1694700623
transform 1 0 196112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_2_2091
timestamp 1694700623
transform 1 0 203952 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1_1326
timestamp 1694700623
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_1_1327
timestamp 1694700623
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2_2092
timestamp 1694700623
transform 1 0 192192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_2_2093
timestamp 1694700623
transform 1 0 200032 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1_1328
timestamp 1694700623
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_1_1329
timestamp 1694700623
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2_2094
timestamp 1694700623
transform 1 0 196112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_2_2095
timestamp 1694700623
transform 1 0 203952 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_1_1330
timestamp 1694700623
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_1_1331
timestamp 1694700623
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_2_2096
timestamp 1694700623
transform 1 0 192192 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_2_2097
timestamp 1694700623
transform 1 0 200032 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_1_1332
timestamp 1694700623
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_1_1333
timestamp 1694700623
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_2_2098
timestamp 1694700623
transform 1 0 196112 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_2_2099
timestamp 1694700623
transform 1 0 203952 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_1_1334
timestamp 1694700623
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_1_1335
timestamp 1694700623
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_2_2100
timestamp 1694700623
transform 1 0 192192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_2_2101
timestamp 1694700623
transform 1 0 200032 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_1_1336
timestamp 1694700623
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_1_1337
timestamp 1694700623
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_2_2102
timestamp 1694700623
transform 1 0 196112 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_2_2103
timestamp 1694700623
transform 1 0 203952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_1_1338
timestamp 1694700623
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_1_1339
timestamp 1694700623
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_2_2104
timestamp 1694700623
transform 1 0 192192 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_2_2105
timestamp 1694700623
transform 1 0 200032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_1_1340
timestamp 1694700623
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_1_1341
timestamp 1694700623
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_2_2106
timestamp 1694700623
transform 1 0 196112 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_2_2107
timestamp 1694700623
transform 1 0 203952 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_1_1342
timestamp 1694700623
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_1_1343
timestamp 1694700623
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_2_2108
timestamp 1694700623
transform 1 0 192192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_2_2109
timestamp 1694700623
transform 1 0 200032 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_1_1344
timestamp 1694700623
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_1_1345
timestamp 1694700623
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_2_2110
timestamp 1694700623
transform 1 0 196112 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_2_2111
timestamp 1694700623
transform 1 0 203952 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_1_1346
timestamp 1694700623
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_1_1347
timestamp 1694700623
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_2_2112
timestamp 1694700623
transform 1 0 192192 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_2_2113
timestamp 1694700623
transform 1 0 200032 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_1_1348
timestamp 1694700623
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_1_1349
timestamp 1694700623
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_2_2114
timestamp 1694700623
transform 1 0 196112 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_2_2115
timestamp 1694700623
transform 1 0 203952 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_1_1350
timestamp 1694700623
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_1_1351
timestamp 1694700623
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_2_2116
timestamp 1694700623
transform 1 0 192192 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_2_2117
timestamp 1694700623
transform 1 0 200032 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_1_1352
timestamp 1694700623
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_1_1353
timestamp 1694700623
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_2_2118
timestamp 1694700623
transform 1 0 196112 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_2_2119
timestamp 1694700623
transform 1 0 203952 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_1_1354
timestamp 1694700623
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_1_1355
timestamp 1694700623
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_2_2120
timestamp 1694700623
transform 1 0 192192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_2_2121
timestamp 1694700623
transform 1 0 200032 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_1_1356
timestamp 1694700623
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_1_1357
timestamp 1694700623
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_2_2122
timestamp 1694700623
transform 1 0 196112 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_2_2123
timestamp 1694700623
transform 1 0 203952 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_1_1358
timestamp 1694700623
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_1_1359
timestamp 1694700623
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_2_2124
timestamp 1694700623
transform 1 0 192192 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_2_2125
timestamp 1694700623
transform 1 0 200032 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_1_1360
timestamp 1694700623
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_1_1361
timestamp 1694700623
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_2_2126
timestamp 1694700623
transform 1 0 196112 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_2_2127
timestamp 1694700623
transform 1 0 203952 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1_1362
timestamp 1694700623
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1_1363
timestamp 1694700623
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_2_2128
timestamp 1694700623
transform 1 0 192192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_2_2129
timestamp 1694700623
transform 1 0 200032 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1_1364
timestamp 1694700623
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1_1365
timestamp 1694700623
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_2_2130
timestamp 1694700623
transform 1 0 196112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_2_2131
timestamp 1694700623
transform 1 0 203952 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1_1366
timestamp 1694700623
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1_1367
timestamp 1694700623
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_2_2132
timestamp 1694700623
transform 1 0 192192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_2_2133
timestamp 1694700623
transform 1 0 200032 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1_1368
timestamp 1694700623
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1_1369
timestamp 1694700623
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_2_2134
timestamp 1694700623
transform 1 0 196112 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_2_2135
timestamp 1694700623
transform 1 0 203952 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1_1370
timestamp 1694700623
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1_1371
timestamp 1694700623
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_2_2136
timestamp 1694700623
transform 1 0 192192 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_2_2137
timestamp 1694700623
transform 1 0 200032 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1_1372
timestamp 1694700623
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1_1373
timestamp 1694700623
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_2_2138
timestamp 1694700623
transform 1 0 196112 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_2_2139
timestamp 1694700623
transform 1 0 203952 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1_1374
timestamp 1694700623
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1_1375
timestamp 1694700623
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_2_2140
timestamp 1694700623
transform 1 0 192192 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_2_2141
timestamp 1694700623
transform 1 0 200032 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1_1376
timestamp 1694700623
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1_1377
timestamp 1694700623
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_2_2142
timestamp 1694700623
transform 1 0 196112 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_2_2143
timestamp 1694700623
transform 1 0 203952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1_1378
timestamp 1694700623
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1_1379
timestamp 1694700623
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_2_2144
timestamp 1694700623
transform 1 0 192192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_2_2145
timestamp 1694700623
transform 1 0 200032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1_1380
timestamp 1694700623
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1_1381
timestamp 1694700623
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_2_2146
timestamp 1694700623
transform 1 0 196112 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_2_2147
timestamp 1694700623
transform 1 0 203952 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_1_1382
timestamp 1694700623
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_1_1383
timestamp 1694700623
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_2_2148
timestamp 1694700623
transform 1 0 192192 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_2_2149
timestamp 1694700623
transform 1 0 200032 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_1_1384
timestamp 1694700623
transform 1 0 9184 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_1_1385
timestamp 1694700623
transform 1 0 17024 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_2_2150
timestamp 1694700623
transform 1 0 196112 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_2_2151
timestamp 1694700623
transform 1 0 203952 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_1_1386
timestamp 1694700623
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_1_1387
timestamp 1694700623
transform 1 0 13104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_2_2152
timestamp 1694700623
transform 1 0 192192 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_2_2153
timestamp 1694700623
transform 1 0 200032 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_1_1388
timestamp 1694700623
transform 1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_1_1389
timestamp 1694700623
transform 1 0 17024 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_2_2154
timestamp 1694700623
transform 1 0 196112 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_2_2155
timestamp 1694700623
transform 1 0 203952 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_1_1390
timestamp 1694700623
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_1_1391
timestamp 1694700623
transform 1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_2_2156
timestamp 1694700623
transform 1 0 192192 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_2_2157
timestamp 1694700623
transform 1 0 200032 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_1_1392
timestamp 1694700623
transform 1 0 9184 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_1_1393
timestamp 1694700623
transform 1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_2_2158
timestamp 1694700623
transform 1 0 196112 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_2_2159
timestamp 1694700623
transform 1 0 203952 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_1_1394
timestamp 1694700623
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_1_1395
timestamp 1694700623
transform 1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_2_2160
timestamp 1694700623
transform 1 0 192192 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_2_2161
timestamp 1694700623
transform 1 0 200032 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_1_1396
timestamp 1694700623
transform 1 0 9184 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_1_1397
timestamp 1694700623
transform 1 0 17024 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_2_2162
timestamp 1694700623
transform 1 0 196112 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_2_2163
timestamp 1694700623
transform 1 0 203952 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_1_1398
timestamp 1694700623
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_1_1399
timestamp 1694700623
transform 1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_2_2164
timestamp 1694700623
transform 1 0 192192 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_2_2165
timestamp 1694700623
transform 1 0 200032 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_1_1400
timestamp 1694700623
transform 1 0 9184 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_1_1401
timestamp 1694700623
transform 1 0 17024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_2_2166
timestamp 1694700623
transform 1 0 196112 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_2_2167
timestamp 1694700623
transform 1 0 203952 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_1_1402
timestamp 1694700623
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_1_1403
timestamp 1694700623
transform 1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_2_2168
timestamp 1694700623
transform 1 0 192192 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_2_2169
timestamp 1694700623
transform 1 0 200032 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_1_1404
timestamp 1694700623
transform 1 0 9184 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_1_1405
timestamp 1694700623
transform 1 0 17024 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_2_2170
timestamp 1694700623
transform 1 0 196112 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_2_2171
timestamp 1694700623
transform 1 0 203952 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_1_1406
timestamp 1694700623
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_1_1407
timestamp 1694700623
transform 1 0 13104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_2_2172
timestamp 1694700623
transform 1 0 192192 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_2_2173
timestamp 1694700623
transform 1 0 200032 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_1_1408
timestamp 1694700623
transform 1 0 9184 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_1_1409
timestamp 1694700623
transform 1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_2_2174
timestamp 1694700623
transform 1 0 196112 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_2_2175
timestamp 1694700623
transform 1 0 203952 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_1_1410
timestamp 1694700623
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_1_1411
timestamp 1694700623
transform 1 0 13104 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_2_2176
timestamp 1694700623
transform 1 0 192192 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_2_2177
timestamp 1694700623
transform 1 0 200032 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_1_1412
timestamp 1694700623
transform 1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_1_1413
timestamp 1694700623
transform 1 0 17024 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_2_2178
timestamp 1694700623
transform 1 0 196112 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_2_2179
timestamp 1694700623
transform 1 0 203952 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_1_1414
timestamp 1694700623
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_1_1415
timestamp 1694700623
transform 1 0 13104 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_2_2180
timestamp 1694700623
transform 1 0 192192 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_2_2181
timestamp 1694700623
transform 1 0 200032 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_1_1416
timestamp 1694700623
transform 1 0 9184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_1_1417
timestamp 1694700623
transform 1 0 17024 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_2_2182
timestamp 1694700623
transform 1 0 196112 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_2_2183
timestamp 1694700623
transform 1 0 203952 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_1_1418
timestamp 1694700623
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_1_1419
timestamp 1694700623
transform 1 0 13104 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_2_2184
timestamp 1694700623
transform 1 0 192192 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_2_2185
timestamp 1694700623
transform 1 0 200032 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_1_1420
timestamp 1694700623
transform 1 0 9184 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_1_1421
timestamp 1694700623
transform 1 0 17024 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_2_2186
timestamp 1694700623
transform 1 0 196112 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_2_2187
timestamp 1694700623
transform 1 0 203952 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_1_1422
timestamp 1694700623
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_1_1423
timestamp 1694700623
transform 1 0 13104 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_2_2188
timestamp 1694700623
transform 1 0 192192 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_2_2189
timestamp 1694700623
transform 1 0 200032 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_1_1424
timestamp 1694700623
transform 1 0 9184 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_1_1425
timestamp 1694700623
transform 1 0 17024 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_2_2190
timestamp 1694700623
transform 1 0 196112 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_2_2191
timestamp 1694700623
transform 1 0 203952 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_1_1426
timestamp 1694700623
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_1_1427
timestamp 1694700623
transform 1 0 13104 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_2_2192
timestamp 1694700623
transform 1 0 192192 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_2_2193
timestamp 1694700623
transform 1 0 200032 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_1_1428
timestamp 1694700623
transform 1 0 9184 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_1_1429
timestamp 1694700623
transform 1 0 17024 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_2_2194
timestamp 1694700623
transform 1 0 196112 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_2_2195
timestamp 1694700623
transform 1 0 203952 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_1_1430
timestamp 1694700623
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_1_1431
timestamp 1694700623
transform 1 0 13104 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_2_2196
timestamp 1694700623
transform 1 0 192192 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_2_2197
timestamp 1694700623
transform 1 0 200032 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_1_1432
timestamp 1694700623
transform 1 0 9184 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_1_1433
timestamp 1694700623
transform 1 0 17024 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_2_2198
timestamp 1694700623
transform 1 0 196112 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_2_2199
timestamp 1694700623
transform 1 0 203952 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_1_1434
timestamp 1694700623
transform 1 0 5264 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_1_1435
timestamp 1694700623
transform 1 0 13104 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_2_2200
timestamp 1694700623
transform 1 0 192192 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_2_2201
timestamp 1694700623
transform 1 0 200032 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_1_1436
timestamp 1694700623
transform 1 0 9184 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_1_1437
timestamp 1694700623
transform 1 0 17024 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_2_2202
timestamp 1694700623
transform 1 0 196112 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_2_2203
timestamp 1694700623
transform 1 0 203952 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_1_1438
timestamp 1694700623
transform 1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_1_1439
timestamp 1694700623
transform 1 0 13104 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_2_2204
timestamp 1694700623
transform 1 0 192192 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_2_2205
timestamp 1694700623
transform 1 0 200032 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_1_1440
timestamp 1694700623
transform 1 0 9184 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_1_1441
timestamp 1694700623
transform 1 0 17024 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_2_2206
timestamp 1694700623
transform 1 0 196112 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_2_2207
timestamp 1694700623
transform 1 0 203952 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_1_1442
timestamp 1694700623
transform 1 0 5264 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_1_1443
timestamp 1694700623
transform 1 0 13104 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_2_2208
timestamp 1694700623
transform 1 0 192192 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_2_2209
timestamp 1694700623
transform 1 0 200032 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_1_1444
timestamp 1694700623
transform 1 0 9184 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_1_1445
timestamp 1694700623
transform 1 0 17024 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_2_2210
timestamp 1694700623
transform 1 0 196112 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_2_2211
timestamp 1694700623
transform 1 0 203952 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_1_1446
timestamp 1694700623
transform 1 0 5264 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_1_1447
timestamp 1694700623
transform 1 0 13104 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_2_2212
timestamp 1694700623
transform 1 0 192192 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_2_2213
timestamp 1694700623
transform 1 0 200032 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_1_1448
timestamp 1694700623
transform 1 0 9184 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_1_1449
timestamp 1694700623
transform 1 0 17024 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_2_2214
timestamp 1694700623
transform 1 0 196112 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_2_2215
timestamp 1694700623
transform 1 0 203952 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_1_1450
timestamp 1694700623
transform 1 0 5264 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_1_1451
timestamp 1694700623
transform 1 0 13104 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_2_2216
timestamp 1694700623
transform 1 0 192192 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_2_2217
timestamp 1694700623
transform 1 0 200032 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_1_1452
timestamp 1694700623
transform 1 0 9184 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_1_1453
timestamp 1694700623
transform 1 0 17024 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_2_2218
timestamp 1694700623
transform 1 0 196112 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_2_2219
timestamp 1694700623
transform 1 0 203952 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_1_1454
timestamp 1694700623
transform 1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_1_1455
timestamp 1694700623
transform 1 0 13104 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_2_2220
timestamp 1694700623
transform 1 0 192192 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_2_2221
timestamp 1694700623
transform 1 0 200032 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_1_1456
timestamp 1694700623
transform 1 0 9184 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_1_1457
timestamp 1694700623
transform 1 0 17024 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_2_2222
timestamp 1694700623
transform 1 0 196112 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_2_2223
timestamp 1694700623
transform 1 0 203952 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_1_1458
timestamp 1694700623
transform 1 0 5264 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_1_1459
timestamp 1694700623
transform 1 0 13104 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_2_2224
timestamp 1694700623
transform 1 0 192192 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_2_2225
timestamp 1694700623
transform 1 0 200032 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_1_1460
timestamp 1694700623
transform 1 0 9184 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_1_1461
timestamp 1694700623
transform 1 0 17024 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_2_2226
timestamp 1694700623
transform 1 0 196112 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_2_2227
timestamp 1694700623
transform 1 0 203952 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_1_1462
timestamp 1694700623
transform 1 0 5264 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_1_1463
timestamp 1694700623
transform 1 0 13104 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_2_2228
timestamp 1694700623
transform 1 0 192192 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_2_2229
timestamp 1694700623
transform 1 0 200032 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_1_1464
timestamp 1694700623
transform 1 0 9184 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_1_1465
timestamp 1694700623
transform 1 0 17024 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_2_2230
timestamp 1694700623
transform 1 0 196112 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_2_2231
timestamp 1694700623
transform 1 0 203952 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_1_1466
timestamp 1694700623
transform 1 0 5264 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_1_1467
timestamp 1694700623
transform 1 0 13104 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_2_2232
timestamp 1694700623
transform 1 0 192192 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_2_2233
timestamp 1694700623
transform 1 0 200032 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_1_1468
timestamp 1694700623
transform 1 0 9184 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_1_1469
timestamp 1694700623
transform 1 0 17024 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_2_2234
timestamp 1694700623
transform 1 0 196112 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_2_2235
timestamp 1694700623
transform 1 0 203952 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_1_1470
timestamp 1694700623
transform 1 0 5264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_1_1471
timestamp 1694700623
transform 1 0 13104 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_2_2236
timestamp 1694700623
transform 1 0 192192 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_2_2237
timestamp 1694700623
transform 1 0 200032 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_1_1472
timestamp 1694700623
transform 1 0 9184 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_1_1473
timestamp 1694700623
transform 1 0 17024 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_2_2238
timestamp 1694700623
transform 1 0 196112 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_2_2239
timestamp 1694700623
transform 1 0 203952 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_1_1474
timestamp 1694700623
transform 1 0 5264 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_1_1475
timestamp 1694700623
transform 1 0 13104 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_2_2240
timestamp 1694700623
transform 1 0 192192 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_2_2241
timestamp 1694700623
transform 1 0 200032 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_1_1476
timestamp 1694700623
transform 1 0 9184 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_1_1477
timestamp 1694700623
transform 1 0 17024 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_2_2242
timestamp 1694700623
transform 1 0 196112 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_2_2243
timestamp 1694700623
transform 1 0 203952 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_1_1478
timestamp 1694700623
transform 1 0 5264 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_1_1479
timestamp 1694700623
transform 1 0 13104 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_2_2244
timestamp 1694700623
transform 1 0 192192 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_2_2245
timestamp 1694700623
transform 1 0 200032 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_1_1480
timestamp 1694700623
transform 1 0 9184 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_1_1481
timestamp 1694700623
transform 1 0 17024 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_2_2246
timestamp 1694700623
transform 1 0 196112 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_2_2247
timestamp 1694700623
transform 1 0 203952 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_1_1482
timestamp 1694700623
transform 1 0 5264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_1_1483
timestamp 1694700623
transform 1 0 13104 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_2_2248
timestamp 1694700623
transform 1 0 192192 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_144_2_2249
timestamp 1694700623
transform 1 0 200032 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_1_1484
timestamp 1694700623
transform 1 0 9184 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_1_1485
timestamp 1694700623
transform 1 0 17024 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_2_2250
timestamp 1694700623
transform 1 0 196112 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_145_2_2251
timestamp 1694700623
transform 1 0 203952 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_1_1486
timestamp 1694700623
transform 1 0 5264 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_1_1487
timestamp 1694700623
transform 1 0 13104 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_2_2252
timestamp 1694700623
transform 1 0 192192 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_146_2_2253
timestamp 1694700623
transform 1 0 200032 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_1_1488
timestamp 1694700623
transform 1 0 9184 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_1_1489
timestamp 1694700623
transform 1 0 17024 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_2_2254
timestamp 1694700623
transform 1 0 196112 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_147_2_2255
timestamp 1694700623
transform 1 0 203952 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_1_1490
timestamp 1694700623
transform 1 0 5264 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_1_1491
timestamp 1694700623
transform 1 0 13104 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_2_2256
timestamp 1694700623
transform 1 0 192192 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_148_2_2257
timestamp 1694700623
transform 1 0 200032 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_149_1_1492
timestamp 1694700623
transform 1 0 9184 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_149_1_1493
timestamp 1694700623
transform 1 0 17024 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_149_2_2258
timestamp 1694700623
transform 1 0 196112 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_149_2_2259
timestamp 1694700623
transform 1 0 203952 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_150_1_1494
timestamp 1694700623
transform 1 0 5264 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_150_1_1495
timestamp 1694700623
transform 1 0 13104 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_150_2_2260
timestamp 1694700623
transform 1 0 192192 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_150_2_2261
timestamp 1694700623
transform 1 0 200032 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_151_1_1496
timestamp 1694700623
transform 1 0 9184 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_151_1_1497
timestamp 1694700623
transform 1 0 17024 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_151_2_2262
timestamp 1694700623
transform 1 0 196112 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_151_2_2263
timestamp 1694700623
transform 1 0 203952 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_152_1_1498
timestamp 1694700623
transform 1 0 5264 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_152_1_1499
timestamp 1694700623
transform 1 0 13104 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_152_2_2264
timestamp 1694700623
transform 1 0 192192 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_152_2_2265
timestamp 1694700623
transform 1 0 200032 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_153_1_1500
timestamp 1694700623
transform 1 0 9184 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_153_1_1501
timestamp 1694700623
transform 1 0 17024 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_153_2_2266
timestamp 1694700623
transform 1 0 196112 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_153_2_2267
timestamp 1694700623
transform 1 0 203952 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_154_1_1502
timestamp 1694700623
transform 1 0 5264 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_154_1_1503
timestamp 1694700623
transform 1 0 13104 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_154_2_2268
timestamp 1694700623
transform 1 0 192192 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_154_2_2269
timestamp 1694700623
transform 1 0 200032 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_155_1_1504
timestamp 1694700623
transform 1 0 9184 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_155_1_1505
timestamp 1694700623
transform 1 0 17024 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_155_2_2270
timestamp 1694700623
transform 1 0 196112 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_155_2_2271
timestamp 1694700623
transform 1 0 203952 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_156_1_1506
timestamp 1694700623
transform 1 0 5264 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_156_1_1507
timestamp 1694700623
transform 1 0 13104 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_156_2_2272
timestamp 1694700623
transform 1 0 192192 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_156_2_2273
timestamp 1694700623
transform 1 0 200032 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_157_1_1508
timestamp 1694700623
transform 1 0 9184 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_157_1_1509
timestamp 1694700623
transform 1 0 17024 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_157_2_2274
timestamp 1694700623
transform 1 0 196112 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_157_2_2275
timestamp 1694700623
transform 1 0 203952 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_158_1_1510
timestamp 1694700623
transform 1 0 5264 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_158_1_1511
timestamp 1694700623
transform 1 0 13104 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_158_2_2276
timestamp 1694700623
transform 1 0 192192 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_158_2_2277
timestamp 1694700623
transform 1 0 200032 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_159_1_1512
timestamp 1694700623
transform 1 0 9184 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_159_1_1513
timestamp 1694700623
transform 1 0 17024 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_159_2_2278
timestamp 1694700623
transform 1 0 196112 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_159_2_2279
timestamp 1694700623
transform 1 0 203952 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_160_1_1514
timestamp 1694700623
transform 1 0 5264 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_160_1_1515
timestamp 1694700623
transform 1 0 13104 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_160_2_2280
timestamp 1694700623
transform 1 0 192192 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_160_2_2281
timestamp 1694700623
transform 1 0 200032 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_161_1_1516
timestamp 1694700623
transform 1 0 9184 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_161_1_1517
timestamp 1694700623
transform 1 0 17024 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_161_2_2282
timestamp 1694700623
transform 1 0 196112 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_161_2_2283
timestamp 1694700623
transform 1 0 203952 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_162_1_1518
timestamp 1694700623
transform 1 0 5264 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_162_1_1519
timestamp 1694700623
transform 1 0 13104 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_162_2_2284
timestamp 1694700623
transform 1 0 192192 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_162_2_2285
timestamp 1694700623
transform 1 0 200032 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_163_1_1520
timestamp 1694700623
transform 1 0 9184 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_163_1_1521
timestamp 1694700623
transform 1 0 17024 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_163_2_2286
timestamp 1694700623
transform 1 0 196112 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_163_2_2287
timestamp 1694700623
transform 1 0 203952 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_164_1_1522
timestamp 1694700623
transform 1 0 5264 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_164_1_1523
timestamp 1694700623
transform 1 0 13104 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_164_2_2288
timestamp 1694700623
transform 1 0 192192 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_164_2_2289
timestamp 1694700623
transform 1 0 200032 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_165_1_1524
timestamp 1694700623
transform 1 0 9184 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_165_1_1525
timestamp 1694700623
transform 1 0 17024 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_165_2_2290
timestamp 1694700623
transform 1 0 196112 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_165_2_2291
timestamp 1694700623
transform 1 0 203952 0 -1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_166_1_1526
timestamp 1694700623
transform 1 0 5264 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_166_1_1527
timestamp 1694700623
transform 1 0 13104 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_166_2_2292
timestamp 1694700623
transform 1 0 192192 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_166_2_2293
timestamp 1694700623
transform 1 0 200032 0 1 133280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_167_1_1528
timestamp 1694700623
transform 1 0 9184 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_167_1_1529
timestamp 1694700623
transform 1 0 17024 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_167_2_2294
timestamp 1694700623
transform 1 0 196112 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_167_2_2295
timestamp 1694700623
transform 1 0 203952 0 -1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_168_1_1530
timestamp 1694700623
transform 1 0 5264 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_168_1_1531
timestamp 1694700623
transform 1 0 13104 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_168_2_2296
timestamp 1694700623
transform 1 0 192192 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_168_2_2297
timestamp 1694700623
transform 1 0 200032 0 1 134848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_169_1_1532
timestamp 1694700623
transform 1 0 9184 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_169_1_1533
timestamp 1694700623
transform 1 0 17024 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_169_2_2298
timestamp 1694700623
transform 1 0 196112 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_169_2_2299
timestamp 1694700623
transform 1 0 203952 0 -1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_170_1_1534
timestamp 1694700623
transform 1 0 5264 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_170_1_1535
timestamp 1694700623
transform 1 0 13104 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_170_2_2300
timestamp 1694700623
transform 1 0 192192 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_170_2_2301
timestamp 1694700623
transform 1 0 200032 0 1 136416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_171_1_1536
timestamp 1694700623
transform 1 0 9184 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_171_1_1537
timestamp 1694700623
transform 1 0 17024 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_171_2_2302
timestamp 1694700623
transform 1 0 196112 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_171_2_2303
timestamp 1694700623
transform 1 0 203952 0 -1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_172_1_1538
timestamp 1694700623
transform 1 0 5264 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_172_1_1539
timestamp 1694700623
transform 1 0 13104 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_172_2_2304
timestamp 1694700623
transform 1 0 192192 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_172_2_2305
timestamp 1694700623
transform 1 0 200032 0 1 137984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_173_1_1540
timestamp 1694700623
transform 1 0 9184 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_173_1_1541
timestamp 1694700623
transform 1 0 17024 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_173_2_2306
timestamp 1694700623
transform 1 0 196112 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_173_2_2307
timestamp 1694700623
transform 1 0 203952 0 -1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_174_1_1542
timestamp 1694700623
transform 1 0 5264 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_174_1_1543
timestamp 1694700623
transform 1 0 13104 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_174_2_2308
timestamp 1694700623
transform 1 0 192192 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_174_2_2309
timestamp 1694700623
transform 1 0 200032 0 1 139552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_175_1_1544
timestamp 1694700623
transform 1 0 9184 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_175_1_1545
timestamp 1694700623
transform 1 0 17024 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_175_2_2310
timestamp 1694700623
transform 1 0 196112 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_175_2_2311
timestamp 1694700623
transform 1 0 203952 0 -1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_176_1_1546
timestamp 1694700623
transform 1 0 5264 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_176_1_1547
timestamp 1694700623
transform 1 0 13104 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_176_2_2312
timestamp 1694700623
transform 1 0 192192 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_176_2_2313
timestamp 1694700623
transform 1 0 200032 0 1 141120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_177_1_1548
timestamp 1694700623
transform 1 0 9184 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_177_1_1549
timestamp 1694700623
transform 1 0 17024 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_177_2_2314
timestamp 1694700623
transform 1 0 196112 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_177_2_2315
timestamp 1694700623
transform 1 0 203952 0 -1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_178_1_1550
timestamp 1694700623
transform 1 0 5264 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_178_1_1551
timestamp 1694700623
transform 1 0 13104 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_178_2_2316
timestamp 1694700623
transform 1 0 192192 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_178_2_2317
timestamp 1694700623
transform 1 0 200032 0 1 142688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_179_1_1552
timestamp 1694700623
transform 1 0 9184 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_179_1_1553
timestamp 1694700623
transform 1 0 17024 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_179_2_2318
timestamp 1694700623
transform 1 0 196112 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_179_2_2319
timestamp 1694700623
transform 1 0 203952 0 -1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_180_1_1554
timestamp 1694700623
transform 1 0 5264 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_180_1_1555
timestamp 1694700623
transform 1 0 13104 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_180_2_2320
timestamp 1694700623
transform 1 0 192192 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_180_2_2321
timestamp 1694700623
transform 1 0 200032 0 1 144256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1556
timestamp 1694700623
transform 1 0 5152 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1557
timestamp 1694700623
transform 1 0 8960 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1558
timestamp 1694700623
transform 1 0 12768 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1559
timestamp 1694700623
transform 1 0 16576 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1560
timestamp 1694700623
transform 1 0 20384 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1561
timestamp 1694700623
transform 1 0 24192 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1562
timestamp 1694700623
transform 1 0 28000 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1563
timestamp 1694700623
transform 1 0 31808 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1564
timestamp 1694700623
transform 1 0 35616 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1565
timestamp 1694700623
transform 1 0 39424 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1566
timestamp 1694700623
transform 1 0 43232 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1567
timestamp 1694700623
transform 1 0 47040 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1568
timestamp 1694700623
transform 1 0 50848 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1569
timestamp 1694700623
transform 1 0 54656 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1570
timestamp 1694700623
transform 1 0 58464 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1571
timestamp 1694700623
transform 1 0 62272 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1572
timestamp 1694700623
transform 1 0 66080 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1573
timestamp 1694700623
transform 1 0 69888 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1574
timestamp 1694700623
transform 1 0 73696 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1575
timestamp 1694700623
transform 1 0 77504 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1576
timestamp 1694700623
transform 1 0 81312 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1577
timestamp 1694700623
transform 1 0 85120 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1578
timestamp 1694700623
transform 1 0 88928 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1579
timestamp 1694700623
transform 1 0 92736 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1580
timestamp 1694700623
transform 1 0 96544 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1581
timestamp 1694700623
transform 1 0 100352 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1582
timestamp 1694700623
transform 1 0 104160 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1583
timestamp 1694700623
transform 1 0 107968 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1584
timestamp 1694700623
transform 1 0 111776 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1585
timestamp 1694700623
transform 1 0 115584 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1586
timestamp 1694700623
transform 1 0 119392 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1587
timestamp 1694700623
transform 1 0 123200 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1588
timestamp 1694700623
transform 1 0 127008 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1589
timestamp 1694700623
transform 1 0 130816 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1590
timestamp 1694700623
transform 1 0 134624 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1591
timestamp 1694700623
transform 1 0 138432 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1592
timestamp 1694700623
transform 1 0 142240 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1593
timestamp 1694700623
transform 1 0 146048 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1594
timestamp 1694700623
transform 1 0 149856 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1595
timestamp 1694700623
transform 1 0 153664 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1596
timestamp 1694700623
transform 1 0 157472 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1597
timestamp 1694700623
transform 1 0 161280 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1598
timestamp 1694700623
transform 1 0 165088 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1599
timestamp 1694700623
transform 1 0 168896 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1600
timestamp 1694700623
transform 1 0 172704 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1601
timestamp 1694700623
transform 1 0 176512 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1602
timestamp 1694700623
transform 1 0 180320 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1603
timestamp 1694700623
transform 1 0 184128 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1604
timestamp 1694700623
transform 1 0 187936 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1605
timestamp 1694700623
transform 1 0 191744 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1606
timestamp 1694700623
transform 1 0 195552 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1607
timestamp 1694700623
transform 1 0 199360 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_181_1608
timestamp 1694700623
transform 1 0 203168 0 -1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1609
timestamp 1694700623
transform 1 0 5264 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1610
timestamp 1694700623
transform 1 0 13104 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1611
timestamp 1694700623
transform 1 0 20944 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1612
timestamp 1694700623
transform 1 0 28784 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1613
timestamp 1694700623
transform 1 0 36624 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1614
timestamp 1694700623
transform 1 0 44464 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1615
timestamp 1694700623
transform 1 0 52304 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1616
timestamp 1694700623
transform 1 0 60144 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1617
timestamp 1694700623
transform 1 0 67984 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1618
timestamp 1694700623
transform 1 0 75824 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1619
timestamp 1694700623
transform 1 0 83664 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1620
timestamp 1694700623
transform 1 0 91504 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1621
timestamp 1694700623
transform 1 0 99344 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1622
timestamp 1694700623
transform 1 0 107184 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1623
timestamp 1694700623
transform 1 0 115024 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1624
timestamp 1694700623
transform 1 0 122864 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1625
timestamp 1694700623
transform 1 0 130704 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1626
timestamp 1694700623
transform 1 0 138544 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1627
timestamp 1694700623
transform 1 0 146384 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1628
timestamp 1694700623
transform 1 0 154224 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1629
timestamp 1694700623
transform 1 0 162064 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1630
timestamp 1694700623
transform 1 0 169904 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1631
timestamp 1694700623
transform 1 0 177744 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1632
timestamp 1694700623
transform 1 0 185584 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1633
timestamp 1694700623
transform 1 0 193424 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_182_1634
timestamp 1694700623
transform 1 0 201264 0 1 145824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1635
timestamp 1694700623
transform 1 0 9184 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1636
timestamp 1694700623
transform 1 0 17024 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1637
timestamp 1694700623
transform 1 0 24864 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1638
timestamp 1694700623
transform 1 0 32704 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1639
timestamp 1694700623
transform 1 0 40544 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1640
timestamp 1694700623
transform 1 0 48384 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1641
timestamp 1694700623
transform 1 0 56224 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1642
timestamp 1694700623
transform 1 0 64064 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1643
timestamp 1694700623
transform 1 0 71904 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1644
timestamp 1694700623
transform 1 0 79744 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1645
timestamp 1694700623
transform 1 0 87584 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1646
timestamp 1694700623
transform 1 0 95424 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1647
timestamp 1694700623
transform 1 0 103264 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1648
timestamp 1694700623
transform 1 0 111104 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1649
timestamp 1694700623
transform 1 0 118944 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1650
timestamp 1694700623
transform 1 0 126784 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1651
timestamp 1694700623
transform 1 0 134624 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1652
timestamp 1694700623
transform 1 0 142464 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1653
timestamp 1694700623
transform 1 0 150304 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1654
timestamp 1694700623
transform 1 0 158144 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1655
timestamp 1694700623
transform 1 0 165984 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1656
timestamp 1694700623
transform 1 0 173824 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1657
timestamp 1694700623
transform 1 0 181664 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1658
timestamp 1694700623
transform 1 0 189504 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_183_1659
timestamp 1694700623
transform 1 0 197344 0 -1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1660
timestamp 1694700623
transform 1 0 5264 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1661
timestamp 1694700623
transform 1 0 13104 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1662
timestamp 1694700623
transform 1 0 20944 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1663
timestamp 1694700623
transform 1 0 28784 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1664
timestamp 1694700623
transform 1 0 36624 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1665
timestamp 1694700623
transform 1 0 44464 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1666
timestamp 1694700623
transform 1 0 52304 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1667
timestamp 1694700623
transform 1 0 60144 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1668
timestamp 1694700623
transform 1 0 67984 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1669
timestamp 1694700623
transform 1 0 75824 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1670
timestamp 1694700623
transform 1 0 83664 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1671
timestamp 1694700623
transform 1 0 91504 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1672
timestamp 1694700623
transform 1 0 99344 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1673
timestamp 1694700623
transform 1 0 107184 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1674
timestamp 1694700623
transform 1 0 115024 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1675
timestamp 1694700623
transform 1 0 122864 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1676
timestamp 1694700623
transform 1 0 130704 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1677
timestamp 1694700623
transform 1 0 138544 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1678
timestamp 1694700623
transform 1 0 146384 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1679
timestamp 1694700623
transform 1 0 154224 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1680
timestamp 1694700623
transform 1 0 162064 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1681
timestamp 1694700623
transform 1 0 169904 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1682
timestamp 1694700623
transform 1 0 177744 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1683
timestamp 1694700623
transform 1 0 185584 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1684
timestamp 1694700623
transform 1 0 193424 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_184_1685
timestamp 1694700623
transform 1 0 201264 0 1 147392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1686
timestamp 1694700623
transform 1 0 9184 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1687
timestamp 1694700623
transform 1 0 17024 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1688
timestamp 1694700623
transform 1 0 24864 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1689
timestamp 1694700623
transform 1 0 32704 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1690
timestamp 1694700623
transform 1 0 40544 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1691
timestamp 1694700623
transform 1 0 48384 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1692
timestamp 1694700623
transform 1 0 56224 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1693
timestamp 1694700623
transform 1 0 64064 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1694
timestamp 1694700623
transform 1 0 71904 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1695
timestamp 1694700623
transform 1 0 79744 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1696
timestamp 1694700623
transform 1 0 87584 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1697
timestamp 1694700623
transform 1 0 95424 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1698
timestamp 1694700623
transform 1 0 103264 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1699
timestamp 1694700623
transform 1 0 111104 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1700
timestamp 1694700623
transform 1 0 118944 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1701
timestamp 1694700623
transform 1 0 126784 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1702
timestamp 1694700623
transform 1 0 134624 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1703
timestamp 1694700623
transform 1 0 142464 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1704
timestamp 1694700623
transform 1 0 150304 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1705
timestamp 1694700623
transform 1 0 158144 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1706
timestamp 1694700623
transform 1 0 165984 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1707
timestamp 1694700623
transform 1 0 173824 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1708
timestamp 1694700623
transform 1 0 181664 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1709
timestamp 1694700623
transform 1 0 189504 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_185_1710
timestamp 1694700623
transform 1 0 197344 0 -1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1711
timestamp 1694700623
transform 1 0 5264 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1712
timestamp 1694700623
transform 1 0 13104 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1713
timestamp 1694700623
transform 1 0 20944 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1714
timestamp 1694700623
transform 1 0 28784 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1715
timestamp 1694700623
transform 1 0 36624 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1716
timestamp 1694700623
transform 1 0 44464 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1717
timestamp 1694700623
transform 1 0 52304 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1718
timestamp 1694700623
transform 1 0 60144 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1719
timestamp 1694700623
transform 1 0 67984 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1720
timestamp 1694700623
transform 1 0 75824 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1721
timestamp 1694700623
transform 1 0 83664 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1722
timestamp 1694700623
transform 1 0 91504 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1723
timestamp 1694700623
transform 1 0 99344 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1724
timestamp 1694700623
transform 1 0 107184 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1725
timestamp 1694700623
transform 1 0 115024 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1726
timestamp 1694700623
transform 1 0 122864 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1727
timestamp 1694700623
transform 1 0 130704 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1728
timestamp 1694700623
transform 1 0 138544 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1729
timestamp 1694700623
transform 1 0 146384 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1730
timestamp 1694700623
transform 1 0 154224 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1731
timestamp 1694700623
transform 1 0 162064 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1732
timestamp 1694700623
transform 1 0 169904 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1733
timestamp 1694700623
transform 1 0 177744 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1734
timestamp 1694700623
transform 1 0 185584 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1735
timestamp 1694700623
transform 1 0 193424 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_186_1736
timestamp 1694700623
transform 1 0 201264 0 1 148960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1737
timestamp 1694700623
transform 1 0 9184 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1738
timestamp 1694700623
transform 1 0 17024 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1739
timestamp 1694700623
transform 1 0 24864 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1740
timestamp 1694700623
transform 1 0 32704 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1741
timestamp 1694700623
transform 1 0 40544 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1742
timestamp 1694700623
transform 1 0 48384 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1743
timestamp 1694700623
transform 1 0 56224 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1744
timestamp 1694700623
transform 1 0 64064 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1745
timestamp 1694700623
transform 1 0 71904 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1746
timestamp 1694700623
transform 1 0 79744 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1747
timestamp 1694700623
transform 1 0 87584 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1748
timestamp 1694700623
transform 1 0 95424 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1749
timestamp 1694700623
transform 1 0 103264 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1750
timestamp 1694700623
transform 1 0 111104 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1751
timestamp 1694700623
transform 1 0 118944 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1752
timestamp 1694700623
transform 1 0 126784 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1753
timestamp 1694700623
transform 1 0 134624 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1754
timestamp 1694700623
transform 1 0 142464 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1755
timestamp 1694700623
transform 1 0 150304 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1756
timestamp 1694700623
transform 1 0 158144 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1757
timestamp 1694700623
transform 1 0 165984 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1758
timestamp 1694700623
transform 1 0 173824 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1759
timestamp 1694700623
transform 1 0 181664 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1760
timestamp 1694700623
transform 1 0 189504 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_187_1761
timestamp 1694700623
transform 1 0 197344 0 -1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1762
timestamp 1694700623
transform 1 0 5264 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1763
timestamp 1694700623
transform 1 0 13104 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1764
timestamp 1694700623
transform 1 0 20944 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1765
timestamp 1694700623
transform 1 0 28784 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1766
timestamp 1694700623
transform 1 0 36624 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1767
timestamp 1694700623
transform 1 0 44464 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1768
timestamp 1694700623
transform 1 0 52304 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1769
timestamp 1694700623
transform 1 0 60144 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1770
timestamp 1694700623
transform 1 0 67984 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1771
timestamp 1694700623
transform 1 0 75824 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1772
timestamp 1694700623
transform 1 0 83664 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1773
timestamp 1694700623
transform 1 0 91504 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1774
timestamp 1694700623
transform 1 0 99344 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1775
timestamp 1694700623
transform 1 0 107184 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1776
timestamp 1694700623
transform 1 0 115024 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1777
timestamp 1694700623
transform 1 0 122864 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1778
timestamp 1694700623
transform 1 0 130704 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1779
timestamp 1694700623
transform 1 0 138544 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1780
timestamp 1694700623
transform 1 0 146384 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1781
timestamp 1694700623
transform 1 0 154224 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1782
timestamp 1694700623
transform 1 0 162064 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1783
timestamp 1694700623
transform 1 0 169904 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1784
timestamp 1694700623
transform 1 0 177744 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1785
timestamp 1694700623
transform 1 0 185584 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1786
timestamp 1694700623
transform 1 0 193424 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_188_1787
timestamp 1694700623
transform 1 0 201264 0 1 150528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1788
timestamp 1694700623
transform 1 0 9184 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1789
timestamp 1694700623
transform 1 0 17024 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1790
timestamp 1694700623
transform 1 0 24864 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1791
timestamp 1694700623
transform 1 0 32704 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1792
timestamp 1694700623
transform 1 0 40544 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1793
timestamp 1694700623
transform 1 0 48384 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1794
timestamp 1694700623
transform 1 0 56224 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1795
timestamp 1694700623
transform 1 0 64064 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1796
timestamp 1694700623
transform 1 0 71904 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1797
timestamp 1694700623
transform 1 0 79744 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1798
timestamp 1694700623
transform 1 0 87584 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1799
timestamp 1694700623
transform 1 0 95424 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1800
timestamp 1694700623
transform 1 0 103264 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1801
timestamp 1694700623
transform 1 0 111104 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1802
timestamp 1694700623
transform 1 0 118944 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1803
timestamp 1694700623
transform 1 0 126784 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1804
timestamp 1694700623
transform 1 0 134624 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1805
timestamp 1694700623
transform 1 0 142464 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1806
timestamp 1694700623
transform 1 0 150304 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1807
timestamp 1694700623
transform 1 0 158144 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1808
timestamp 1694700623
transform 1 0 165984 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1809
timestamp 1694700623
transform 1 0 173824 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1810
timestamp 1694700623
transform 1 0 181664 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1811
timestamp 1694700623
transform 1 0 189504 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_189_1812
timestamp 1694700623
transform 1 0 197344 0 -1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1813
timestamp 1694700623
transform 1 0 5264 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1814
timestamp 1694700623
transform 1 0 13104 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1815
timestamp 1694700623
transform 1 0 20944 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1816
timestamp 1694700623
transform 1 0 28784 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1817
timestamp 1694700623
transform 1 0 36624 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1818
timestamp 1694700623
transform 1 0 44464 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1819
timestamp 1694700623
transform 1 0 52304 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1820
timestamp 1694700623
transform 1 0 60144 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1821
timestamp 1694700623
transform 1 0 67984 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1822
timestamp 1694700623
transform 1 0 75824 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1823
timestamp 1694700623
transform 1 0 83664 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1824
timestamp 1694700623
transform 1 0 91504 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1825
timestamp 1694700623
transform 1 0 99344 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1826
timestamp 1694700623
transform 1 0 107184 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1827
timestamp 1694700623
transform 1 0 115024 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1828
timestamp 1694700623
transform 1 0 122864 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1829
timestamp 1694700623
transform 1 0 130704 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1830
timestamp 1694700623
transform 1 0 138544 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1831
timestamp 1694700623
transform 1 0 146384 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1832
timestamp 1694700623
transform 1 0 154224 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1833
timestamp 1694700623
transform 1 0 162064 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1834
timestamp 1694700623
transform 1 0 169904 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1835
timestamp 1694700623
transform 1 0 177744 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1836
timestamp 1694700623
transform 1 0 185584 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1837
timestamp 1694700623
transform 1 0 193424 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_190_1838
timestamp 1694700623
transform 1 0 201264 0 1 152096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1839
timestamp 1694700623
transform 1 0 9184 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1840
timestamp 1694700623
transform 1 0 17024 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1841
timestamp 1694700623
transform 1 0 24864 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1842
timestamp 1694700623
transform 1 0 32704 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1843
timestamp 1694700623
transform 1 0 40544 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1844
timestamp 1694700623
transform 1 0 48384 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1845
timestamp 1694700623
transform 1 0 56224 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1846
timestamp 1694700623
transform 1 0 64064 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1847
timestamp 1694700623
transform 1 0 71904 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1848
timestamp 1694700623
transform 1 0 79744 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1849
timestamp 1694700623
transform 1 0 87584 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1850
timestamp 1694700623
transform 1 0 95424 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1851
timestamp 1694700623
transform 1 0 103264 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1852
timestamp 1694700623
transform 1 0 111104 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1853
timestamp 1694700623
transform 1 0 118944 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1854
timestamp 1694700623
transform 1 0 126784 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1855
timestamp 1694700623
transform 1 0 134624 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1856
timestamp 1694700623
transform 1 0 142464 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1857
timestamp 1694700623
transform 1 0 150304 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1858
timestamp 1694700623
transform 1 0 158144 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1859
timestamp 1694700623
transform 1 0 165984 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1860
timestamp 1694700623
transform 1 0 173824 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1861
timestamp 1694700623
transform 1 0 181664 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1862
timestamp 1694700623
transform 1 0 189504 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_191_1863
timestamp 1694700623
transform 1 0 197344 0 -1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1864
timestamp 1694700623
transform 1 0 5264 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1865
timestamp 1694700623
transform 1 0 13104 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1866
timestamp 1694700623
transform 1 0 20944 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1867
timestamp 1694700623
transform 1 0 28784 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1868
timestamp 1694700623
transform 1 0 36624 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1869
timestamp 1694700623
transform 1 0 44464 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1870
timestamp 1694700623
transform 1 0 52304 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1871
timestamp 1694700623
transform 1 0 60144 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1872
timestamp 1694700623
transform 1 0 67984 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1873
timestamp 1694700623
transform 1 0 75824 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1874
timestamp 1694700623
transform 1 0 83664 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1875
timestamp 1694700623
transform 1 0 91504 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1876
timestamp 1694700623
transform 1 0 99344 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1877
timestamp 1694700623
transform 1 0 107184 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1878
timestamp 1694700623
transform 1 0 115024 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1879
timestamp 1694700623
transform 1 0 122864 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1880
timestamp 1694700623
transform 1 0 130704 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1881
timestamp 1694700623
transform 1 0 138544 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1882
timestamp 1694700623
transform 1 0 146384 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1883
timestamp 1694700623
transform 1 0 154224 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1884
timestamp 1694700623
transform 1 0 162064 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1885
timestamp 1694700623
transform 1 0 169904 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1886
timestamp 1694700623
transform 1 0 177744 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1887
timestamp 1694700623
transform 1 0 185584 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1888
timestamp 1694700623
transform 1 0 193424 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_192_1889
timestamp 1694700623
transform 1 0 201264 0 1 153664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1890
timestamp 1694700623
transform 1 0 9184 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1891
timestamp 1694700623
transform 1 0 17024 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1892
timestamp 1694700623
transform 1 0 24864 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1893
timestamp 1694700623
transform 1 0 32704 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1894
timestamp 1694700623
transform 1 0 40544 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1895
timestamp 1694700623
transform 1 0 48384 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1896
timestamp 1694700623
transform 1 0 56224 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1897
timestamp 1694700623
transform 1 0 64064 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1898
timestamp 1694700623
transform 1 0 71904 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1899
timestamp 1694700623
transform 1 0 79744 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1900
timestamp 1694700623
transform 1 0 87584 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1901
timestamp 1694700623
transform 1 0 95424 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1902
timestamp 1694700623
transform 1 0 103264 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1903
timestamp 1694700623
transform 1 0 111104 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1904
timestamp 1694700623
transform 1 0 118944 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1905
timestamp 1694700623
transform 1 0 126784 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1906
timestamp 1694700623
transform 1 0 134624 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1907
timestamp 1694700623
transform 1 0 142464 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1908
timestamp 1694700623
transform 1 0 150304 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1909
timestamp 1694700623
transform 1 0 158144 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1910
timestamp 1694700623
transform 1 0 165984 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1911
timestamp 1694700623
transform 1 0 173824 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1912
timestamp 1694700623
transform 1 0 181664 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1913
timestamp 1694700623
transform 1 0 189504 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_193_1914
timestamp 1694700623
transform 1 0 197344 0 -1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1915
timestamp 1694700623
transform 1 0 5264 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1916
timestamp 1694700623
transform 1 0 13104 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1917
timestamp 1694700623
transform 1 0 20944 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1918
timestamp 1694700623
transform 1 0 28784 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1919
timestamp 1694700623
transform 1 0 36624 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1920
timestamp 1694700623
transform 1 0 44464 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1921
timestamp 1694700623
transform 1 0 52304 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1922
timestamp 1694700623
transform 1 0 60144 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1923
timestamp 1694700623
transform 1 0 67984 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1924
timestamp 1694700623
transform 1 0 75824 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1925
timestamp 1694700623
transform 1 0 83664 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1926
timestamp 1694700623
transform 1 0 91504 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1927
timestamp 1694700623
transform 1 0 99344 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1928
timestamp 1694700623
transform 1 0 107184 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1929
timestamp 1694700623
transform 1 0 115024 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1930
timestamp 1694700623
transform 1 0 122864 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1931
timestamp 1694700623
transform 1 0 130704 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1932
timestamp 1694700623
transform 1 0 138544 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1933
timestamp 1694700623
transform 1 0 146384 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1934
timestamp 1694700623
transform 1 0 154224 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1935
timestamp 1694700623
transform 1 0 162064 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1936
timestamp 1694700623
transform 1 0 169904 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1937
timestamp 1694700623
transform 1 0 177744 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1938
timestamp 1694700623
transform 1 0 185584 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1939
timestamp 1694700623
transform 1 0 193424 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_194_1940
timestamp 1694700623
transform 1 0 201264 0 1 155232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1941
timestamp 1694700623
transform 1 0 5152 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1942
timestamp 1694700623
transform 1 0 8960 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1943
timestamp 1694700623
transform 1 0 12768 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1944
timestamp 1694700623
transform 1 0 16576 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1945
timestamp 1694700623
transform 1 0 20384 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1946
timestamp 1694700623
transform 1 0 24192 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1947
timestamp 1694700623
transform 1 0 28000 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1948
timestamp 1694700623
transform 1 0 31808 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1949
timestamp 1694700623
transform 1 0 35616 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1950
timestamp 1694700623
transform 1 0 39424 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1951
timestamp 1694700623
transform 1 0 43232 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1952
timestamp 1694700623
transform 1 0 47040 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1953
timestamp 1694700623
transform 1 0 50848 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1954
timestamp 1694700623
transform 1 0 54656 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1955
timestamp 1694700623
transform 1 0 58464 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1956
timestamp 1694700623
transform 1 0 62272 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1957
timestamp 1694700623
transform 1 0 66080 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1958
timestamp 1694700623
transform 1 0 69888 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1959
timestamp 1694700623
transform 1 0 73696 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1960
timestamp 1694700623
transform 1 0 77504 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1961
timestamp 1694700623
transform 1 0 81312 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1962
timestamp 1694700623
transform 1 0 85120 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1963
timestamp 1694700623
transform 1 0 88928 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1964
timestamp 1694700623
transform 1 0 92736 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1965
timestamp 1694700623
transform 1 0 96544 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1966
timestamp 1694700623
transform 1 0 100352 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1967
timestamp 1694700623
transform 1 0 104160 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1968
timestamp 1694700623
transform 1 0 107968 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1969
timestamp 1694700623
transform 1 0 111776 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1970
timestamp 1694700623
transform 1 0 115584 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1971
timestamp 1694700623
transform 1 0 119392 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1972
timestamp 1694700623
transform 1 0 123200 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1973
timestamp 1694700623
transform 1 0 127008 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1974
timestamp 1694700623
transform 1 0 130816 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1975
timestamp 1694700623
transform 1 0 134624 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1976
timestamp 1694700623
transform 1 0 138432 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1977
timestamp 1694700623
transform 1 0 142240 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1978
timestamp 1694700623
transform 1 0 146048 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1979
timestamp 1694700623
transform 1 0 149856 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1980
timestamp 1694700623
transform 1 0 153664 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1981
timestamp 1694700623
transform 1 0 157472 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1982
timestamp 1694700623
transform 1 0 161280 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1983
timestamp 1694700623
transform 1 0 165088 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1984
timestamp 1694700623
transform 1 0 168896 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1985
timestamp 1694700623
transform 1 0 172704 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1986
timestamp 1694700623
transform 1 0 176512 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1987
timestamp 1694700623
transform 1 0 180320 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1988
timestamp 1694700623
transform 1 0 184128 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1989
timestamp 1694700623
transform 1 0 187936 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1990
timestamp 1694700623
transform 1 0 191744 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1991
timestamp 1694700623
transform 1 0 195552 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1992
timestamp 1694700623
transform 1 0 199360 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_195_1993
timestamp 1694700623
transform 1 0 203168 0 -1 156800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_30 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 149072 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_31
timestamp 1694700623
transform -1 0 126224 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_32
timestamp 1694700623
transform -1 0 103376 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_33
timestamp 1694700623
transform -1 0 80528 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_34
timestamp 1694700623
transform -1 0 57680 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_35
timestamp 1694700623
transform -1 0 34832 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_36
timestamp 1694700623
transform -1 0 11984 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_37
timestamp 1694700623
transform -1 0 2016 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_38
timestamp 1694700623
transform -1 0 2016 0 1 142688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_39
timestamp 1694700623
transform -1 0 2016 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_40
timestamp 1694700623
transform -1 0 2016 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_41
timestamp 1694700623
transform -1 0 2016 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_42
timestamp 1694700623
transform -1 0 2016 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_43
timestamp 1694700623
transform -1 0 2016 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_44
timestamp 1694700623
transform -1 0 2016 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_45
timestamp 1694700623
transform -1 0 2016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_46
timestamp 1694700623
transform -1 0 2016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_47
timestamp 1694700623
transform -1 0 2016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_48
timestamp 1694700623
transform -1 0 2016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_49
timestamp 1694700623
transform -1 0 2016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_50
timestamp 1694700623
transform -1 0 2016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_51
timestamp 1694700623
transform -1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_52
timestamp 1694700623
transform -1 0 103376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_53
timestamp 1694700623
transform -1 0 171920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_54
timestamp 1694700623
transform 1 0 204064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_55
timestamp 1694700623
transform 1 0 203504 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_56
timestamp 1694700623
transform 1 0 204064 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_57
timestamp 1694700623
transform 1 0 204064 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_58
timestamp 1694700623
transform 1 0 203504 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_59
timestamp 1694700623
transform 1 0 204064 0 -1 155232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_60
timestamp 1694700623
transform -1 0 187152 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  user_proj_example_61
timestamp 1694700623
transform -1 0 164304 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_62 pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 95760 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_63
timestamp 1694700623
transform -1 0 72912 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_64
timestamp 1694700623
transform -1 0 50064 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_65
timestamp 1694700623
transform -1 0 27216 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_66
timestamp 1694700623
transform -1 0 4368 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_67
timestamp 1694700623
transform -1 0 2016 0 1 150528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_68
timestamp 1694700623
transform -1 0 2016 0 -1 139552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_69
timestamp 1694700623
transform -1 0 2016 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_70
timestamp 1694700623
transform -1 0 2016 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_71
timestamp 1694700623
transform -1 0 2016 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_72
timestamp 1694700623
transform -1 0 2016 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_73
timestamp 1694700623
transform -1 0 2016 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_74
timestamp 1694700623
transform -1 0 2016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_75
timestamp 1694700623
transform -1 0 2016 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_76
timestamp 1694700623
transform -1 0 2016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_77
timestamp 1694700623
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_78
timestamp 1694700623
transform -1 0 2016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_79
timestamp 1694700623
transform -1 0 2016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_80
timestamp 1694700623
transform -1 0 2016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_81
timestamp 1694700623
transform -1 0 141456 0 -1 156800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  user_proj_example_82
timestamp 1694700623
transform -1 0 118608 0 -1 156800
box -86 -86 534 870
<< labels >>
flabel metal3 s 205332 5600 206132 5712 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 110432 159264 110544 160064 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 87584 159264 87696 160064 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 64736 159264 64848 160064 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 41888 159264 42000 160064 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 19040 159264 19152 160064 0 FreeSans 448 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal3 s 0 157920 800 158032 0 FreeSans 448 0 0 0 io_in[15]
port 6 nsew signal input
flabel metal3 s 0 146496 800 146608 0 FreeSans 448 0 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 0 135072 800 135184 0 FreeSans 448 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal3 s 0 123648 800 123760 0 FreeSans 448 0 0 0 io_in[18]
port 9 nsew signal input
flabel metal3 s 0 112224 800 112336 0 FreeSans 448 0 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 205332 31808 206132 31920 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal3 s 0 100800 800 100912 0 FreeSans 448 0 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 0 89376 800 89488 0 FreeSans 448 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal3 s 0 77952 800 78064 0 FreeSans 448 0 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 0 66528 800 66640 0 FreeSans 448 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 55104 800 55216 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 9408 800 9520 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 205332 58016 206132 58128 0 FreeSans 448 0 0 0 io_in[2]
port 21 nsew signal input
flabel metal3 s 205332 84224 206132 84336 0 FreeSans 448 0 0 0 io_in[3]
port 22 nsew signal input
flabel metal3 s 205332 110432 206132 110544 0 FreeSans 448 0 0 0 io_in[4]
port 23 nsew signal input
flabel metal3 s 205332 136640 206132 136752 0 FreeSans 448 0 0 0 io_in[5]
port 24 nsew signal input
flabel metal2 s 201824 159264 201936 160064 0 FreeSans 448 90 0 0 io_in[6]
port 25 nsew signal input
flabel metal2 s 178976 159264 179088 160064 0 FreeSans 448 90 0 0 io_in[7]
port 26 nsew signal input
flabel metal2 s 156128 159264 156240 160064 0 FreeSans 448 90 0 0 io_in[8]
port 27 nsew signal input
flabel metal2 s 133280 159264 133392 160064 0 FreeSans 448 90 0 0 io_in[9]
port 28 nsew signal input
flabel metal3 s 205332 23072 206132 23184 0 FreeSans 448 0 0 0 io_oeb[0]
port 29 nsew signal tristate
flabel metal2 s 95200 159264 95312 160064 0 FreeSans 448 90 0 0 io_oeb[10]
port 30 nsew signal tristate
flabel metal2 s 72352 159264 72464 160064 0 FreeSans 448 90 0 0 io_oeb[11]
port 31 nsew signal tristate
flabel metal2 s 49504 159264 49616 160064 0 FreeSans 448 90 0 0 io_oeb[12]
port 32 nsew signal tristate
flabel metal2 s 26656 159264 26768 160064 0 FreeSans 448 90 0 0 io_oeb[13]
port 33 nsew signal tristate
flabel metal2 s 3808 159264 3920 160064 0 FreeSans 448 90 0 0 io_oeb[14]
port 34 nsew signal tristate
flabel metal3 s 0 150304 800 150416 0 FreeSans 448 0 0 0 io_oeb[15]
port 35 nsew signal tristate
flabel metal3 s 0 138880 800 138992 0 FreeSans 448 0 0 0 io_oeb[16]
port 36 nsew signal tristate
flabel metal3 s 0 127456 800 127568 0 FreeSans 448 0 0 0 io_oeb[17]
port 37 nsew signal tristate
flabel metal3 s 0 116032 800 116144 0 FreeSans 448 0 0 0 io_oeb[18]
port 38 nsew signal tristate
flabel metal3 s 0 104608 800 104720 0 FreeSans 448 0 0 0 io_oeb[19]
port 39 nsew signal tristate
flabel metal3 s 205332 49280 206132 49392 0 FreeSans 448 0 0 0 io_oeb[1]
port 40 nsew signal tristate
flabel metal3 s 0 93184 800 93296 0 FreeSans 448 0 0 0 io_oeb[20]
port 41 nsew signal tristate
flabel metal3 s 0 81760 800 81872 0 FreeSans 448 0 0 0 io_oeb[21]
port 42 nsew signal tristate
flabel metal3 s 0 70336 800 70448 0 FreeSans 448 0 0 0 io_oeb[22]
port 43 nsew signal tristate
flabel metal3 s 0 58912 800 59024 0 FreeSans 448 0 0 0 io_oeb[23]
port 44 nsew signal tristate
flabel metal3 s 0 47488 800 47600 0 FreeSans 448 0 0 0 io_oeb[24]
port 45 nsew signal tristate
flabel metal3 s 0 36064 800 36176 0 FreeSans 448 0 0 0 io_oeb[25]
port 46 nsew signal tristate
flabel metal3 s 0 24640 800 24752 0 FreeSans 448 0 0 0 io_oeb[26]
port 47 nsew signal tristate
flabel metal3 s 0 13216 800 13328 0 FreeSans 448 0 0 0 io_oeb[27]
port 48 nsew signal tristate
flabel metal3 s 0 1792 800 1904 0 FreeSans 448 0 0 0 io_oeb[28]
port 49 nsew signal tristate
flabel metal3 s 205332 75488 206132 75600 0 FreeSans 448 0 0 0 io_oeb[2]
port 50 nsew signal tristate
flabel metal3 s 205332 101696 206132 101808 0 FreeSans 448 0 0 0 io_oeb[3]
port 51 nsew signal tristate
flabel metal3 s 205332 127904 206132 128016 0 FreeSans 448 0 0 0 io_oeb[4]
port 52 nsew signal tristate
flabel metal3 s 205332 154112 206132 154224 0 FreeSans 448 0 0 0 io_oeb[5]
port 53 nsew signal tristate
flabel metal2 s 186592 159264 186704 160064 0 FreeSans 448 90 0 0 io_oeb[6]
port 54 nsew signal tristate
flabel metal2 s 163744 159264 163856 160064 0 FreeSans 448 90 0 0 io_oeb[7]
port 55 nsew signal tristate
flabel metal2 s 140896 159264 141008 160064 0 FreeSans 448 90 0 0 io_oeb[8]
port 56 nsew signal tristate
flabel metal2 s 118048 159264 118160 160064 0 FreeSans 448 90 0 0 io_oeb[9]
port 57 nsew signal tristate
flabel metal3 s 205332 14336 206132 14448 0 FreeSans 448 0 0 0 io_out[0]
port 58 nsew signal tristate
flabel metal2 s 102816 159264 102928 160064 0 FreeSans 448 90 0 0 io_out[10]
port 59 nsew signal tristate
flabel metal2 s 79968 159264 80080 160064 0 FreeSans 448 90 0 0 io_out[11]
port 60 nsew signal tristate
flabel metal2 s 57120 159264 57232 160064 0 FreeSans 448 90 0 0 io_out[12]
port 61 nsew signal tristate
flabel metal2 s 34272 159264 34384 160064 0 FreeSans 448 90 0 0 io_out[13]
port 62 nsew signal tristate
flabel metal2 s 11424 159264 11536 160064 0 FreeSans 448 90 0 0 io_out[14]
port 63 nsew signal tristate
flabel metal3 s 0 154112 800 154224 0 FreeSans 448 0 0 0 io_out[15]
port 64 nsew signal tristate
flabel metal3 s 0 142688 800 142800 0 FreeSans 448 0 0 0 io_out[16]
port 65 nsew signal tristate
flabel metal3 s 0 131264 800 131376 0 FreeSans 448 0 0 0 io_out[17]
port 66 nsew signal tristate
flabel metal3 s 0 119840 800 119952 0 FreeSans 448 0 0 0 io_out[18]
port 67 nsew signal tristate
flabel metal3 s 0 108416 800 108528 0 FreeSans 448 0 0 0 io_out[19]
port 68 nsew signal tristate
flabel metal3 s 205332 40544 206132 40656 0 FreeSans 448 0 0 0 io_out[1]
port 69 nsew signal tristate
flabel metal3 s 0 96992 800 97104 0 FreeSans 448 0 0 0 io_out[20]
port 70 nsew signal tristate
flabel metal3 s 0 85568 800 85680 0 FreeSans 448 0 0 0 io_out[21]
port 71 nsew signal tristate
flabel metal3 s 0 74144 800 74256 0 FreeSans 448 0 0 0 io_out[22]
port 72 nsew signal tristate
flabel metal3 s 0 62720 800 62832 0 FreeSans 448 0 0 0 io_out[23]
port 73 nsew signal tristate
flabel metal3 s 0 51296 800 51408 0 FreeSans 448 0 0 0 io_out[24]
port 74 nsew signal tristate
flabel metal3 s 0 39872 800 39984 0 FreeSans 448 0 0 0 io_out[25]
port 75 nsew signal tristate
flabel metal3 s 0 28448 800 28560 0 FreeSans 448 0 0 0 io_out[26]
port 76 nsew signal tristate
flabel metal3 s 0 17024 800 17136 0 FreeSans 448 0 0 0 io_out[27]
port 77 nsew signal tristate
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 io_out[28]
port 78 nsew signal tristate
flabel metal3 s 205332 66752 206132 66864 0 FreeSans 448 0 0 0 io_out[2]
port 79 nsew signal tristate
flabel metal3 s 205332 92960 206132 93072 0 FreeSans 448 0 0 0 io_out[3]
port 80 nsew signal tristate
flabel metal3 s 205332 119168 206132 119280 0 FreeSans 448 0 0 0 io_out[4]
port 81 nsew signal tristate
flabel metal3 s 205332 145376 206132 145488 0 FreeSans 448 0 0 0 io_out[5]
port 82 nsew signal tristate
flabel metal2 s 194208 159264 194320 160064 0 FreeSans 448 90 0 0 io_out[6]
port 83 nsew signal tristate
flabel metal2 s 171360 159264 171472 160064 0 FreeSans 448 90 0 0 io_out[7]
port 84 nsew signal tristate
flabel metal2 s 148512 159264 148624 160064 0 FreeSans 448 90 0 0 io_out[8]
port 85 nsew signal tristate
flabel metal2 s 125664 159264 125776 160064 0 FreeSans 448 90 0 0 io_out[9]
port 86 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 irq[0]
port 87 nsew signal tristate
flabel metal2 s 102816 0 102928 800 0 FreeSans 448 90 0 0 irq[1]
port 88 nsew signal tristate
flabel metal2 s 171360 0 171472 800 0 FreeSans 448 90 0 0 irq[2]
port 89 nsew signal tristate
flabel metal4 s 4448 3076 4768 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 35168 3076 35488 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 65888 3076 66208 20065 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 65888 142955 66208 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 96608 3076 96928 17888 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 96608 39876 96928 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 127328 3076 127648 21188 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 127328 35384 127648 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 158048 3076 158368 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 188768 3076 189088 156860 0 FreeSans 1280 90 0 0 vdd
port 90 nsew power bidirectional
flabel metal5 s 1284 6306 204796 6626 0 FreeSans 2304 0 0 0 vdd
port 90 nsew power bidirectional
flabel metal5 s 1284 36942 204796 37262 0 FreeSans 2304 0 0 0 vdd
port 90 nsew power bidirectional
flabel metal5 s 1284 67578 204796 67898 0 FreeSans 2304 0 0 0 vdd
port 90 nsew power bidirectional
flabel metal5 s 1284 98214 204796 98534 0 FreeSans 2304 0 0 0 vdd
port 90 nsew power bidirectional
flabel metal5 s 1284 128850 204796 129170 0 FreeSans 2304 0 0 0 vdd
port 90 nsew power bidirectional
flabel metal4 s 5108 3076 5428 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 35828 3076 36148 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 66548 3076 66868 20065 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 66548 35384 66868 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 97268 3076 97588 21056 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 97268 35384 97588 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 127988 3076 128308 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 158708 3076 159028 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal4 s 189428 3076 189748 156860 0 FreeSans 1280 90 0 0 vss
port 91 nsew ground bidirectional
flabel metal5 s 1284 6966 204796 7286 0 FreeSans 2304 0 0 0 vss
port 91 nsew ground bidirectional
flabel metal5 s 1284 37602 204796 37922 0 FreeSans 2304 0 0 0 vss
port 91 nsew ground bidirectional
flabel metal5 s 1284 68238 204796 68558 0 FreeSans 2304 0 0 0 vss
port 91 nsew ground bidirectional
flabel metal5 s 1284 98874 204796 99194 0 FreeSans 2304 0 0 0 vss
port 91 nsew ground bidirectional
flabel metal5 s 1284 129510 204796 129830 0 FreeSans 2304 0 0 0 vss
port 91 nsew ground bidirectional
rlabel via4 185538 129114 185538 129114 0 vdd
rlabel via4 186198 129774 186198 129774 0 vss
rlabel metal2 110488 157962 110488 157962 0 io_in[10]
rlabel metal2 88536 156744 88536 156744 0 io_in[11]
rlabel metal2 64792 157850 64792 157850 0 io_in[12]
rlabel metal2 41944 157850 41944 157850 0 io_in[13]
rlabel metal2 19096 157962 19096 157962 0 io_in[14]
rlabel metal2 1736 157192 1736 157192 0 io_in[15]
rlabel metal2 1848 146440 1848 146440 0 io_in[16]
rlabel metal2 1736 135184 1736 135184 0 io_in[17]
rlabel metal3 1302 123704 1302 123704 0 io_in[18]
rlabel metal2 1736 112392 1736 112392 0 io_in[19]
rlabel metal2 1736 101192 1736 101192 0 io_in[20]
rlabel metal2 1736 89488 1736 89488 0 io_in[21]
rlabel metal2 1736 78288 1736 78288 0 io_in[22]
rlabel metal2 1736 66808 1736 66808 0 io_in[23]
rlabel metal3 1246 55160 1246 55160 0 io_in[24]
rlabel metal3 1302 43736 1302 43736 0 io_in[25]
rlabel metal2 1736 32424 1736 32424 0 io_in[26]
rlabel metal2 1736 21224 1736 21224 0 io_in[27]
rlabel metal2 1736 9520 1736 9520 0 io_in[28]
rlabel metal2 157080 156744 157080 156744 0 io_in[8]
rlabel metal2 134232 156912 134232 156912 0 io_in[9]
rlabel metal2 204120 14504 204120 14504 0 io_out[0]
rlabel metal2 204120 40936 204120 40936 0 io_out[1]
rlabel metal2 203224 66864 203224 66864 0 io_out[2]
rlabel metal2 203224 93296 203224 93296 0 io_out[3]
rlabel metal2 204120 119504 204120 119504 0 io_out[4]
rlabel metal2 204120 145880 204120 145880 0 io_out[5]
rlabel metal2 194936 155792 194936 155792 0 io_out[6]
rlabel metal2 171864 156632 171864 156632 0 io_out[7]
rlabel metal3 65240 22246 65240 22246 0 net1
rlabel metal4 54683 21690 54683 21690 0 net10
rlabel metal3 4816 101640 4816 101640 0 net11
rlabel metal2 2184 76860 2184 76860 0 net12
rlabel metal2 2072 77112 2072 77112 0 net13
rlabel metal2 2296 71764 2296 71764 0 net14
rlabel metal3 9128 55272 9128 55272 0 net15
rlabel metal3 8288 44296 8288 44296 0 net16
rlabel metal2 2072 34496 2072 34496 0 net17
rlabel metal2 2128 21784 2128 21784 0 net18
rlabel metal3 7392 9576 7392 9576 0 net19
rlabel metal4 68547 21690 68547 21690 0 net2
rlabel metal4 156408 46368 156408 46368 0 net20
rlabel metal3 61768 22246 61768 22246 0 net21
rlabel via3 67816 20435 67816 20435 0 net22
rlabel metal4 78680 23240 78680 23240 0 net23
rlabel metal2 78904 24080 78904 24080 0 net24
rlabel metal4 77224 23240 77224 23240 0 net25
rlabel via3 125384 26025 125384 26025 0 net26
rlabel via3 140056 26171 140056 26171 0 net27
rlabel metal3 154448 20440 154448 20440 0 net28
rlabel metal2 174048 43848 174048 43848 0 net29
rlabel metal3 72072 22246 72072 22246 0 net3
rlabel metal2 148680 156632 148680 156632 0 net30
rlabel metal2 125832 156632 125832 156632 0 net31
rlabel metal2 102984 156632 102984 156632 0 net32
rlabel metal2 80136 156632 80136 156632 0 net33
rlabel metal2 57288 156632 57288 156632 0 net34
rlabel metal2 34440 156632 34440 156632 0 net35
rlabel metal2 11592 156632 11592 156632 0 net36
rlabel metal3 1246 154168 1246 154168 0 net37
rlabel metal3 1246 142744 1246 142744 0 net38
rlabel metal3 1246 131320 1246 131320 0 net39
rlabel metal4 75385 21690 75385 21690 0 net4
rlabel metal3 1246 119896 1246 119896 0 net40
rlabel metal3 1246 108472 1246 108472 0 net41
rlabel metal3 1246 97048 1246 97048 0 net42
rlabel metal3 1246 85624 1246 85624 0 net43
rlabel metal3 1246 74200 1246 74200 0 net44
rlabel metal3 1246 62776 1246 62776 0 net45
rlabel metal3 1246 51352 1246 51352 0 net46
rlabel metal3 1246 39928 1246 39928 0 net47
rlabel metal3 1246 28504 1246 28504 0 net48
rlabel metal3 1246 17080 1246 17080 0 net49
rlabel metal2 22792 87360 22792 87360 0 net5
rlabel metal3 1246 5656 1246 5656 0 net50
rlabel metal2 34328 2030 34328 2030 0 net51
rlabel metal2 102872 2030 102872 2030 0 net52
rlabel metal2 171416 2030 171416 2030 0 net53
rlabel metal2 204344 23408 204344 23408 0 net54
rlabel metal2 203784 49616 203784 49616 0 net55
rlabel metal3 204890 75544 204890 75544 0 net56
rlabel metal2 204344 101920 204344 101920 0 net57
rlabel metal2 203784 128128 203784 128128 0 net58
rlabel metal2 204344 154560 204344 154560 0 net59
rlabel metal2 75656 24920 75656 24920 0 net6
rlabel metal2 186760 156632 186760 156632 0 net60
rlabel metal2 163912 156632 163912 156632 0 net61
rlabel metal2 95368 156184 95368 156184 0 net62
rlabel metal2 72520 156184 72520 156184 0 net63
rlabel metal2 49672 156184 49672 156184 0 net64
rlabel metal2 26824 156184 26824 156184 0 net65
rlabel metal2 3976 156184 3976 156184 0 net66
rlabel metal3 1246 150360 1246 150360 0 net67
rlabel metal3 1246 138936 1246 138936 0 net68
rlabel metal3 1246 127512 1246 127512 0 net69
rlabel metal4 44373 21690 44373 21690 0 net7
rlabel metal3 1246 116088 1246 116088 0 net70
rlabel metal3 1246 104664 1246 104664 0 net71
rlabel metal3 1246 93240 1246 93240 0 net72
rlabel metal3 1246 81816 1246 81816 0 net73
rlabel metal3 1246 70392 1246 70392 0 net74
rlabel metal3 1246 58968 1246 58968 0 net75
rlabel metal3 1246 47544 1246 47544 0 net76
rlabel metal3 1246 36120 1246 36120 0 net77
rlabel metal3 1246 24696 1246 24696 0 net78
rlabel metal3 1246 13272 1246 13272 0 net79
rlabel via3 48328 20435 48328 20435 0 net8
rlabel metal3 1246 1848 1246 1848 0 net80
rlabel metal2 141064 156184 141064 156184 0 net81
rlabel metal2 118216 156184 118216 156184 0 net82
rlabel metal3 51464 22246 51464 22246 0 net9
<< properties >>
string FIXED_BBOX 0 0 206132 160064
<< end >>
